// See LICENSE.TT for license details.
// Open Vector Interface wrapper module for Ocelot
module tt_vpu_ovi #(parameter VLEN = 256)
(                 input  logic clk, reset_n,

                  input  logic [31:0] issue_inst,
                  input  logic [4:0]  issue_sb_id,
                  input  logic [63:0] issue_scalar_opnd,
                  input  logic [39:0] issue_vcsr,
                  input  logic        issue_vcsr_lmulb2, // Added 1 more bit for vlmul
                  input  logic        issue_valid,
                  output logic        issue_credit,

                  input  logic [4:0]  dispatch_sb_id,
                  input  logic        dispatch_next_senior,
                  input  logic        dispatch_kill,

                  output logic        completed_valid,
                  output logic [4:0]  completed_sb_id,
                  output logic [4:0]  completed_fflags,
                  output logic [63:0] completed_dest_reg,
                  output logic        completed_vxsat,
                  output logic [13:0] completed_vstart,
                  output logic        completed_illegal,

                  output logic         store_valid,
                  output logic [511:0] store_data,
                  input  logic         store_credit,

                  input  logic [33:0]  load_seq_id,
                  input  logic [511:0] load_data,
                  input  logic         load_valid,
                  input  logic [63:0]  load_mask,
                  input  logic         load_mask_valid,

                  input  logic         memop_sync_end,
                  output logic         memop_sync_start,

                  // Debug signals for cosim checker
                  output logic              debug_wb_vec_valid,
                  output logic [VLEN*8-1:0] debug_wb_vec_wdata,
                  output logic [7:0]        debug_wb_vec_wmask
);
                  // TODO: Add the signals for memory operations...

  localparam LOCAL_MEM_BYTE_ADDR_WIDTH = 12;
  localparam INCL_VEC = 1;
//  localparam VLEN = 256;
  localparam ADDRWIDTH = 48;
  localparam LD_DATA_WIDTH_BITS = VLEN;
  localparam ST_DATA_WIDTH_BITS = VLEN;
  localparam LQ_DEPTH=8;
  localparam LQ_DEPTH_LOG2=$clog2(LQ_DEPTH);
  localparam DATA_REQ_ID_WIDTH=INCL_VEC ? (LQ_DEPTH_LOG2+$clog2(VLEN/8)+2) : LQ_DEPTH_LOG2;
  localparam INCL_FP = 1;
  localparam STORE_CREDITS = 32;

  localparam                                          FLEN    = 32;
  localparam                                          FP_RF_RD_PORTS  = 4;
  localparam                                          FP_RF_WR_PORTS  = 2;
  localparam                                          FP_RF_ADDR_WIDTH    = 5;
  localparam                                          EXP_WIDTH   = 8;
  localparam                                          MAN_WIDTH   = 23;
  localparam                                          RS1_IDX = 0;
  localparam                                          RS2_IDX = 1;
  localparam                                          RS3_IDX = 2;

  /////////
  // MEM signals
  wire                     mem_dst_vld;  // forwarding control to ID
  wire [LQ_DEPTH_LOG2-1:0] mem_dst_lqid; // forwarding control to ID
  wire [31:0]              mem_fwd_data; // forwarding control to ID
  wire                     mem_ex_rtr           ;
  wire [ 6:0]              mem_lq_op            ; // mem status to ID
  wire                     mem_lq_commit        ;
    
  tt_briscv_pkg::arr_lq_info_s  lq_broadside_info;
  logic [LQ_DEPTH-1:0][31:0]    lq_broadside_data;
  logic [LQ_DEPTH-1:0]          lq_broadside_valid;
  logic [LQ_DEPTH-1:0]          lq_broadside_data_valid;
  logic                         lq_empty;

  /////////
  // ID signals
  wire                             id_rtr               ;
  wire [4:0]                       id_type              ;
  wire                             id_rf_wr_flag        ;
  wire [ 4:0]                      id_rf_wraddr         ;
  wire                             id_fp_rf_wr_flag     ;
  wire [ 4:0]                      id_fp_rf_wraddr      ;
  wire [31:0]                      id_immed_op          ;
  wire                             id_ex_rts            ;
  wire                             id_ex_units_rts      ;
  wire [LQ_DEPTH_LOG2-1:0]         id_ex_lqid;
  wire [4:0]                       id_ex_Zb_instr       ;
  wire                             id_ex_vecldst        ;
  wire [VLEN-1:0]                  vmask_rddata        ;
  wire [VLEN-1:0]                  vs2_rddata          ; 
  wire [VLEN-1:0]                  vs3_rddata          ; 
  wire [31:0]                      id_ex_pc             ;
  wire                             id_vex_rts           ;
  wire                             vex_id_rtr           ;
  wire [31:0]                      id_ex_instrn         ;
  wire                             v_vm                 ;
  logic [4:0]                      iterate_addrp0,iterate_addrp1,iterate_addrp2       ;
  logic                            ignore_lmul,ignore_dstincr,ignore_srcincr;
  wire [3:0]                       id_fp_fmt             ;
  tt_briscv_pkg::vec_autogen_s     id_vec_autogen;
  tt_briscv_pkg::vecldst_autogen_s id_ex_vecldst_autogen;
  wire                             id_ex_instdisp       ;

  logic                     id_replay;              // From id of tt_id.v
  logic [LQ_DEPTH_LOG2-1:0] id_vex_lqid;          // From id of tt_id.v
  logic                     vex_id_incr_addrp2;     // From vecu of tt_vec.v

  logic                           i_rd_data_vld_2      ;
  logic [DATA_REQ_ID_WIDTH-1:0]   i_rd_data_resp_id_2  ; 

  // Vector signals
  logic              vrf_p0_rden, vrf_p1_rden, vrf_p2_rden;
  logic [VLEN  -1:0] vrf_vm0_rddata;
  logic [VLEN  -1:0] vrf_p0_rddata, vrf_p1_rddata, vrf_p2_rddata;
  logic [       4:0] vrf_p0_rdaddr, vrf_p1_rdaddr, vrf_p2_rdaddr;
  logic              mem_rf_wr;
  logic [       4:0] mem_rf_wraddr;
  logic [      63:0] mem_rf_wrdata;
  logic              mem_fp_rf_wr;
  logic [       4:0] mem_fp_rf_wraddr;
  logic [      63:0] mem_fp_rf_wrdata;
  logic              mem_vrf_wr;
  logic [       4:0] mem_vrf_wraddr;
  logic [VLEN  -1:0] mem_vrf_wrdata;
  logic [VLEN*8-1:0] mem_vrf_wrdata_reg;
  logic [VLEN*8-1:0] mem_vrf_wrdata_nxt;
  logic [       4:0] mem_vrf_wrexc;
  logic [       4:0] mem_vrf_wrexc_reg;
  logic [       4:0] mem_vrf_wrexc_nxt;
  logic [       7:0] mem_vrf_wrmask_reg;
  logic [       7:0] mem_vrf_wrmask_nxt;
  
  logic         vec_store_commit;
  logic         vec_nonstore_commit;

  // LQ signals
  // ID <--> MEM signals
  logic                     mem_fe_lqfull;
  logic                     mem_fe_lqempty;
  logic                     mem_fe_skidbuffull;
  logic [LQ_DEPTH_LOG2-1:0] mem_id_lqnxtid;
  logic [LQ_DEPTH_LOG2-1:0] mem_id_lqnxtid_r;
  logic                     id_mem_lqalloc;
  logic                     id_mem_lq_done;
  tt_briscv_pkg::lq_info_s  id_mem_lqinfo;
  
  // EX --> ID signals
  wire                     ex_dst_vld_1c;
  wire [LQ_DEPTH_LOG2-1:0] ex_dst_lqid_1c;
  wire [31:0]              ex_fwd_data_1c;
    
  wire                     ex_dst_vld_2c;
  wire [LQ_DEPTH_LOG2-1:0] ex_dst_lqid_2c;
  wire [31:0]              ex_fwd_data_2c;
  wire                     ex_id_rtr;
  
  // EX --> MEM signals
  tt_briscv_pkg::mem_skidbuf_s ex_mem_payload;
  wire                         ex_mem_vld           ;

  logic                        ex_mem_lqvld_1c;
  logic [31:0]                 ex_mem_lqdata_1c;
  logic [LQ_DEPTH_LOG2-1:0]    ex_mem_lqid_1c;
    
  logic                        ex_mem_lqvld_2c;
  logic [31:0]                 ex_mem_lqdata_2c;
  logic [LQ_DEPTH_LOG2-1:0]    ex_mem_lqid_2c;
    
  // VEX --> MEM signals
  logic                     vex_mem_lqvld_1c;
  logic [VLEN-1:0]          vex_mem_lqdata_1c;
  logic [LQ_DEPTH_LOG2-1:0] vex_mem_lqid_1c;
  tt_briscv_pkg::csr_fp_exc vex_mem_lqexc_1c;
                        
  logic                     vex_mem_lqvld_2c;
  logic [VLEN-1:0]          vex_mem_lqdata_2c;
  logic [LQ_DEPTH_LOG2-1:0] vex_mem_lqid_2c;
  tt_briscv_pkg::csr_fp_exc vex_mem_lqexc_2c;
                        
  logic                     vex_mem_lqvld_3c;
  logic [VLEN-1:0]          vex_mem_lqdata_3c;
  logic [LQ_DEPTH_LOG2-1:0] vex_mem_lqid_3c;
  tt_briscv_pkg::csr_fp_exc vex_mem_lqexc_3c;

  logic [63:0]  rf_vex_p0_reg;
  logic [63:0]  rf_vex_p1_reg;
  logic [63:0]  fprf_vex_p0_reg;

  logic [63:0]  rf_vex_p0_sel;
  logic [63:0]  rf_vex_p1_sel;
  logic [63:0]  fprf_vex_p0_sel;

 // stall the ID stage when there is a load/store 
  logic ovi_stall;
  logic ocelot_read_req;

  logic        read_valid;
  logic [31:0] read_issue_inst;
  logic [4:0]  read_issue_sb_id;
  logic [63:0] read_issue_scalar_opnd;
  logic [39:0] read_issue_vcsr;
  logic        read_issue_vcsr_lmulb2;

  // I'm using dummy wires to connect the memory interface for now
  logic o_data_req;
  logic [ADDRWIDTH-1:0] o_data_addr;
  logic [ST_DATA_WIDTH_BITS/8-1:0] o_data_byten;
  logic [ST_DATA_WIDTH_BITS-1:0] o_wr_data;
  logic [DATA_REQ_ID_WIDTH-1:0] o_data_req_id;
  logic o_mem_load;
  logic [2:0] o_mem_size;
  logic o_mem_last;

  logic [VLEN*8-1:0] ocelot_instrn_commit_data;
  logic [7:0] ocelot_instrn_commit_mask;
  logic [4:0] ocelot_instrn_commit_fflags;
  logic       ocelot_sat_csr;
  logic       ocelot_instrn_commit_valid;

  // Hack to keep the vector CSRs constant for ocelot
  logic [39:0] vcsr_reg;
  logic        vcsr_lmulb2_reg;
  logic [39:0] vcsr;
  logic        vcsr_lmulb2;

  // Store logic
  logic [7:0][VLEN-1:0] store_buffer;
  logic [7:0] store_buffer_valid;
  // Indicates if the corresponding entry was sent to the CPU
  logic [7:0] store_buffer_sent;
  logic [2:0] store_buffer_wptr;
  logic [2:0] store_buffer_rptr;
  logic [1:0] store_fsm_state; // 0: idle, 1: busy, 2: commit
  logic [1:0] store_fsm_next_state;
  logic       store_memsync_start;
  logic [$clog2(STORE_CREDITS):0] store_credits;
  logic       vecldst_autogen_store;
  // Indicates if there is at least 2 full entries in the store buffer
  logic       enough_data;
  logic       store_buffer_full;
  // This will drive completed.valid
  logic       store_commit;
  // Load logic - finite state machine
  logic [1:0] load_fsm_state, load_fsm_next_state;
  logic       vecldst_autogen_load;
  logic       load_commit;
  logic       load_memsync_start;

  logic [VLEN-1:0][DATA_REQ_ID_WIDTH-1:0] req_buffer;
  logic [$clog2(VLEN)-1:0] req_buffer_wptr;

  logic [511:0] packed_load_data;
  logic [511:0] shifted_load_data;
  logic [4:0]   v_reg;
  logic [10:0]  el_id;
  logic [5:0]   el_off;
  logic [6:0]   el_count;
  logic [4:0]   sb_id;
  // from 0 to 3, 8-bit to 64-bit EEW
  logic [1:0]   eew;
  logic [2:0]   eew_log2;
  // this is in bytes
  logic [63:0]  load_stride;
  // this is in EEW(1,2,4)
  logic [2:0]   load_stride_in_eew_log2;
  // this is the offset of the first element in the packed load data
  logic [5:0] packed_offset;
  logic [10:0] offset_diff;
  logic [$clog2(VLEN)-1:0] shamt;
  logic [8:0] el_id_lower_bound;
  logic [8:0] el_id_upper_bound;
  logic [7:0][VLEN-1:0] load_buffer;  

  always_ff @(posedge clk) begin
    if(!reset_n) begin
      rf_vex_p0_reg   <= '0;
      rf_vex_p1_reg   <= '0;
      fprf_vex_p0_reg <= '0;
    end
    else if (read_valid &&
        ocelot_read_req   ) begin
        rf_vex_p0_reg   <= read_issue_scalar_opnd;
        rf_vex_p1_reg   <= read_issue_scalar_opnd;
        fprf_vex_p0_reg <= read_issue_scalar_opnd;
    end
  end

  assign rf_vex_p0_sel   = (read_valid && ocelot_read_req) ? read_issue_scalar_opnd   : rf_vex_p0_reg;
  assign rf_vex_p1_sel   = (read_valid && ocelot_read_req) ? read_issue_scalar_opnd   : rf_vex_p1_reg;
  assign fprf_vex_p0_sel = (read_valid && ocelot_read_req) ? read_issue_scalar_opnd : fprf_vex_p0_reg;

  tt_briscv_pkg::csr_to_id ex_id_csr;
  assign ex_id_csr.vgsrc   = 0;
  assign ex_id_csr.v_vsew  = vcsr[38:36];
  assign ex_id_csr.v_lmul  = {vcsr_lmulb2,vcsr[35:34]};
  assign ex_id_csr.v_vlmax = '0;
  assign ex_id_csr.v_vl    = vcsr[$clog2(VLEN+1)-1+14:14];

  tt_id
  #(
    .LQ_DEPTH(LQ_DEPTH),
    .LQ_DEPTH_LOG2(LQ_DEPTH_LOG2), 
    .EXP_WIDTH(EXP_WIDTH),
    .MAN_WIDTH(MAN_WIDTH),
    .FLEN(FLEN),
    .VLEN(VLEN),
    .FP_RF_RD_PORTS(FP_RF_RD_PORTS),
    .INCL_VEC(INCL_VEC),
    .INCL_FP(INCL_FP)
  ) id
  (
    .i_clk                                 (clk             ),    
    .i_reset_n                             (reset_n), 

    .i_ex_id_csr                           (ex_id_csr),             

    .i_if_instrn                           (read_issue_inst),       
    .i_if_pc                               ('0),           
    .i_if_instrn_rts                       (read_valid),    
    .o_id_instrn_rtr                       (ocelot_read_req),    

    .o_id_type                             (id_type),          
    .o_id_immed_op                         (id_immed_op),     

    // Vector Interface
    .o_id_vex_rts                          (id_vex_rts),            
    .i_vex_id_rtr                          (vex_id_rtr),            
    .o_vec_autogen                         (id_vec_autogen),   
    .o_id_vex_lqid                         (id_vex_lqid), 
    .i_vex_id_incr_addrp2                  (vex_id_incr_addrp2),    
    .o_v_vm                                (v_vm              ),    

    // EX Interface
    .o_id_ex_rts                           (id_ex_rts),             
    .i_ex_rtr                              (ex_id_rtr         ),    
    .o_id_ex_pc                            (id_ex_pc),        
    .o_id_ex_instrn                        (id_ex_instrn),    
    .o_id_ex_lqid                          (id_ex_lqid[LQ_DEPTH_LOG2-1:0]), 
    .o_id_ex_vecldst                       (id_ex_vecldst),         
    .o_id_ex_Zb_instr                      (id_ex_Zb_instr[4:0]),   
    .o_id_ex_units_rts                     (id_ex_units_rts),       
    .o_id_ex_instdisp                      (id_ex_instdisp),
    .o_vecldst_autogen                     (id_ex_vecldst_autogen), 
    .i_ex_bp_mispredict                    ('0),      
    .i_ex_dst_vld_1c                       (ex_dst_vld_1c),         
    .i_ex_dst_lqid_1c                      (ex_dst_lqid_1c), 
    .i_ex_fwd_data_1c                      (ex_fwd_data_1c),  
    .i_ex_dst_vld_2c                       (ex_dst_vld_2c),         
    .i_ex_dst_lqid_2c                      (ex_dst_lqid_2c), 
    .i_ex_fwd_data_2c                      (ex_fwd_data_2c),  
    .o_fwd_p0_reg                          (),      
    .o_fwd_p1_reg                          (),      

    // FP Interface
    .o_id_fp_ex0_rts                       (),         
    .i_fp_ex0_id_rtr                       (1'b1),         
    .o_id_fp_ex0_lqid                      (), 
    .o_ex_autogen                          (),    
    .o_fp_autogen                          (),   
    .o_fp_fwd_sign_reg                     (),     
    .o_fp_fwd_zero_reg                     (),     
    .o_fp_fwd_nan_reg                      (),      
    .o_fp_fwd_inf_reg                      (),      
    .o_fp_fwd_exp_reg                      (),      
    .o_fp_fwd_man_reg                      (),      
    .o_fp_rf_p3_reg                        (),          
    .i_fp_ex_dst_vld_1c                    ('0),      
    .i_fp_ex_dst_lqid_1c                   ('0), 
    .i_fp_ex_fwd_data_1c                   ('0), 
    .i_fp_ex_dst_vld_2c                    ('0),      
    .i_fp_ex_dst_lqid_2c                   ('0), 
    .i_fp_ex_fwd_data_2c                   ('0), 

    // Integer RegFile Interface
    .o_rf_p0_rden                          (),    
    .o_rf_p0_rdaddr                        (),    
    .o_rf_p1_rden                          (),    
    .o_rf_p1_rdaddr                        (),    
    .o_rf_p2_rden                          (),    
    .o_rf_p2_rdaddr                        (),    
    .o_rf_wr_flag                          (id_rf_wr_flag     ),    
    .o_rf_wraddr                           (id_rf_wraddr      ),    

    // FP RegFile Interface
    .i_fp_rf_rd_ret_reg                    ('0),      
    .i_fp_rf_sign                          ('0),     
    .i_fp_rf_zero                          ('0),     
    .i_fp_rf_nan                           ('0),      
    .i_fp_rf_inf                           ('0),      
    .i_fp_rf_exp                           ('0),      
    .i_fp_rf_man                           ('0),      
    .i_rf_p0_reg                           ('0),       
    .i_rf_p1_reg                           ('0),       
    .o_fp_rf_wr_flag                       (id_fp_rf_wr_flag  ),    
    .o_fp_rf_wraddr                        (id_fp_rf_wraddr   ),    

    // Mem Interface
    .i_lq_broadside_info                   (lq_broadside_info),     
    .o_id_mem_lqinfo                       (id_mem_lqinfo),         
    .o_id_replay                           (id_replay),             
    .o_id_mem_lqalloc                      (id_mem_lqalloc),        
    .o_id_mem_lq_done                      (id_mem_lq_done),        
    .i_mem_dst_vld                         (mem_dst_vld          ), 
    .i_mem_dst_lqid                        (mem_dst_lqid         ), 
    .i_mem_fwd_data                        (mem_fwd_data         ), 
    .i_mem_lq_op                           (mem_lq_op[6:0]),        
    .i_mem_lq_commit                       (mem_lq_commit),         
    .i_lq_broadside_data                   (lq_broadside_data),     
    .i_lq_broadside_valid                  (lq_broadside_valid), 
    .i_lq_broadside_data_valid             (lq_broadside_data_valid), 

    // Misc
    .i_iterate_addrp0                      (iterate_addrp0),   
    .i_iterate_addrp1                      (iterate_addrp1),   
    .i_iterate_addrp2                      (iterate_addrp2),   
    .i_ignore_lmul                         (ignore_lmul),           
    .i_ignore_dstincr                      (ignore_dstincr),        
    .i_ignore_srcincr                      (ignore_srcincr),        
    .i_mem_fe_lqfull                       (mem_fe_lqfull),         
    .i_mem_fe_lqempty                      (mem_fe_lqempty),
    .i_mem_fe_skidbuffull                  (mem_fe_skidbuffull),    
    .i_mem_id_lqnxtid                      (mem_id_lqnxtid[LQ_DEPTH_LOG2-1:0]),

    .i_ovi_stall                           (ovi_stall)
  );  

  //////////
  // EX
  tt_briscv_pkg::csr_to_vec ex_vec_csr;
  assign ex_vec_csr.v_vsew =  vcsr[38:36];
  assign ex_vec_csr.v_lmul =  {vcsr_lmulb2,vcsr[35:34]};
  assign ex_vec_csr.v_vxrm =  vcsr[30:29];
  assign ex_vec_csr.v_vl   =  vcsr[$clog2(VLEN+1)-1+14:14];
  assign vecldst_autogen_store = id_ex_vecldst_autogen.store;
  assign vecldst_autogen_load = id_ex_vecldst_autogen.load;

  tt_ex
  #(.INCL_VEC(INCL_VEC),
    .VLEN(VLEN),
    .LQ_DEPTH_LOG2(LQ_DEPTH_LOG2)
  ) ex
  (
    .i_clk               (clk             ),
    .i_reset_n           (reset_n),
    .i_sat_csr           ('0),
    .i_ex_vec_csr        (ex_vec_csr),             
    // From ID
    .i_if_ex_deco        ('0    ),
    .i_if_ex_predicted   ('0    ),
    .i_if_ex_nextinstr   ('0    ),
    .i_exc_fp_ex_update  ('0    ),
    .i_exc_vfp_update    ('0    ),
    
    // From ID
    .i_id_ex_rts         (id_ex_rts         ),
    .o_ex_id_rtr         (ex_id_rtr         ),
    .i_id_type           (id_type           ),
    .i_id_rf_wr_flag     (id_rf_wr_flag     ),
    .i_id_rf_wraddr      (id_rf_wraddr      ),
    .i_id_fp_rf_wr_flag  (id_fp_rf_wr_flag  ),
    .i_id_fp_rf_wraddr   (id_fp_rf_wraddr   ),
    .i_id_immed_op       (id_immed_op       ),
    .i_id_ex_lqid        (id_ex_lqid        ),
    .i_id_ex_pc          (id_ex_pc          ),
    .i_id_ex_instrn      (id_ex_instrn      ),
    .i_id_ex_vecldst     (id_ex_vecldst     ),
    .i_id_ex_Zb_instr    (id_ex_Zb_instr    ),
    .i_id_ex_units_rts   (id_ex_units_rts   ),
    .i_id_ex_instdisp    (id_ex_instdisp    ),
    
    .i_id_ex_vecldst_autogen(id_ex_vecldst_autogen),
    
    // From RF
    .i_rf_p0_reg         (rf_vex_p0_reg),
    .i_rf_p1_reg         (rf_vex_p1_reg),
    .i_fp_rf_p3_reg      ('0),
    
    // From VRF
    .i_vmask_rddata      (vmask_rddata      ),
    .i_vs2_rddata        (vs2_rddata        ),
    .i_vs3_rddata        (vs3_rddata        ),
    
    // From MEM
    .i_mem_ex_rtr        (mem_ex_rtr        ),
    
    // To ID and IF
    .o_ex_bp_fifo_pop    (),
    .o_ex_is_some_branch (),
    .o_ex_branch_taken   (),
    
    .o_ex_bp_mispredict         (),
    .o_ex_bp_mispredict_not_br  (),
    .o_ex_bp_pc                 (),
    .o_ex_id_csr                (),
    .o_ex_vec_csr               (),
    
    .o_ex_dst_vld_1c        (ex_dst_vld_1c        ),
    .o_ex_dst_lqid_1c       (ex_dst_lqid_1c       ),
    .o_ex_fwd_data_1c       (ex_fwd_data_1c       ),
    .o_ex_dst_vld_2c        (ex_dst_vld_2c        ),
    .o_ex_dst_lqid_2c       (ex_dst_lqid_2c       ),
    .o_ex_fwd_data_2c       (ex_fwd_data_2c       ),
    
    // To MEM
    .o_ex_mem_lqvld_1c      (ex_mem_lqvld_1c     ),
    .o_ex_mem_lqid_1c       (ex_mem_lqid_1c      ),
    .o_ex_mem_lqdata_1c     (ex_mem_lqdata_1c    ),
    
    .o_ex_mem_lqvld_2c      (ex_mem_lqvld_2c     ),
    .o_ex_mem_lqid_2c       (ex_mem_lqid_2c      ),
    .o_ex_mem_lqdata_2c     (ex_mem_lqdata_2c    ),
    
    .o_ex_mem_payload       (ex_mem_payload      ),
    .o_ex_mem_vld           (ex_mem_vld          ),
    
    // Debug
    .i_reset_pc             ('0),

    .i_ovi_stall(ovi_stall)
  );

  assign vrf_p2_rden    = id_vec_autogen.rf_rden2; // FIXME | ex_vec_csr.v_lmul[2];
  assign vrf_p1_rden    = id_vec_autogen.rf_rden1;
  assign vrf_p0_rden    = id_vec_autogen.rf_rden0;

  // VRF read data for EX (V-LD/ST)
  assign vmask_rddata  = vrf_vm0_rddata;
  assign vs2_rddata    = vrf_p1_rddata;
  assign vs3_rddata    = vrf_p2_rddata;

  assign vrf_p0_rdaddr =                                  id_vec_autogen.rf_addrp0;
  assign vrf_p1_rdaddr = id_vec_autogen.rf_rd_p2_is_rs2 ? id_vec_autogen.rf_addrp2
                                                        : id_vec_autogen.rf_addrp1;
  assign vrf_p2_rdaddr = id_vec_autogen.rf_rd_p2_is_rs2 ? id_vec_autogen.rf_addrp1
                                                        : id_vec_autogen.rf_addrp2;

  tt_vec_regfile #(.VLEN(VLEN))
  regfile
  (
    .i_clk               (clk),
    .i_reset_n           (reset_n),
    // Outputs
    .o_rddata_0a         ({vrf_p2_rddata,vrf_p1_rddata,vrf_p0_rddata}),
    .o_dstmask_0a        (),
    .o_vm0_0a            (vrf_vm0_rddata),
    // Inputs
    .i_rden_0a           ({vrf_p2_rden,vrf_p1_rden,vrf_p0_rden}),
    .i_wren_0a           (mem_vrf_wr),
    .i_rdaddr_0a         ({vrf_p2_rdaddr, vrf_p1_rdaddr, vrf_p0_rdaddr}),
    .i_wraddr_0a         (mem_vrf_wraddr),
    .i_wrdata_0a         (mem_vrf_wrdata)
  );

  tt_vec #(.VLEN(VLEN),
          .XLEN(64  ) )
  vecu
  (
    .i_clk                 (clk),                 
    .i_reset_n             (reset_n), 
    .i_ex_vec_csr          (ex_vec_csr),             
    .i_csr_frm             (vcsr[33:31]),
    .i_v_vm                (v_vm),                  
    .i_id_vec_autogen      (id_vec_autogen),        
    .o_sat_csr             (ocelot_sat_csr),
    // ID Interface
    .i_id_vex_rts          (id_vex_rts),            
    .o_vex_id_rtr          (vex_id_rtr),            
    .i_id_ex_vecldst       (id_ex_vecldst),         
    .i_id_ex_instrn        (id_ex_instrn),    
    .i_id_replay           (id_replay),             
    .i_id_type             (id_type),          
    .o_vex_id_incr_addrp2  (vex_id_incr_addrp2),    
    .o_iterate_addrp0      (iterate_addrp0),   
    .o_iterate_addrp1      (iterate_addrp1),   
    .o_iterate_addrp2      (iterate_addrp2),   
    .o_ignore_lmul         (ignore_lmul),           
    .o_ignore_dstincr      (ignore_dstincr),        
    .o_ignore_srcincr      (ignore_srcincr),        
    // RegFile Interface
    .i_rf_vex_p0           (rf_vex_p0_sel),       
    .i_fprf_vex_p0         (fprf_vex_p0_sel),
    .i_vrf_p0_rddata       (vrf_p0_rddata),  
    .i_vrf_p1_rddata       (vrf_p1_rddata),  
    .i_vrf_p2_rddata       (vrf_p2_rddata),  
    .i_vrf_vm0_rddata      (vrf_vm0_rddata),
    // Mem Interface
    .o_vex_mem_lqvld_1c    (vex_mem_lqvld_1c),      
    .o_vex_mem_lqdata_1c   (vex_mem_lqdata_1c), 
    .o_vex_mem_lqexc_1c    (vex_mem_lqexc_1c),      
    .o_vex_mem_lqid_1c     (vex_mem_lqid_1c), 
    .o_vex_mem_lqvld_2c    (vex_mem_lqvld_2c),      
    .o_vex_mem_lqdata_2c   (vex_mem_lqdata_2c), 
    .o_vex_mem_lqexc_2c    (vex_mem_lqexc_2c),      
    .o_vex_mem_lqid_2c     (vex_mem_lqid_2c), 
    .o_vex_mem_lqvld_3c    (vex_mem_lqvld_3c),      
    .o_vex_mem_lqdata_3c   (vex_mem_lqdata_3c), 
    .o_vex_mem_lqexc_3c    (vex_mem_lqexc_3c),      
    .o_vex_mem_lqid_3c     (vex_mem_lqid_3c), 
    .i_mem_vrf_wr          (mem_vrf_wr),            
    .i_mem_vrf_wraddr      (mem_vrf_wraddr),   
    .i_mem_vrf_wrdata      (mem_vrf_wrdata), 
    .i_mem_ex_rtr          (mem_ex_rtr)            
  );    

  logic                        o_data_128b          ;  // 128b read (This signal is valid only for reads)
  logic                        o_data_ordered       ;
  logic [ 3:0]                 o_data_reqtype       ;
  logic                           o_data_req_prequal;
  logic                           i_dmem_brisc_memory_idle; 
  logic                           o_mem_store;
  logic                        o_mem_last_raw;

  tt_mem 
  #(
    .LQ_DEPTH(LQ_DEPTH), 
    .LQ_DEPTH_LOG2(LQ_DEPTH_LOG2),
    .VLEN(VLEN),
    .ADDRWIDTH(ADDRWIDTH),
    .LD_DATA_WIDTH_BITS(LD_DATA_WIDTH_BITS),
    .ST_DATA_WIDTH_BITS(ST_DATA_WIDTH_BITS),  
    .LOCAL_MEM_BYTE_ADDR_WIDTH(LOCAL_MEM_BYTE_ADDR_WIDTH),
    .DATA_REQ_ID_WIDTH(DATA_REQ_ID_WIDTH),
    .INCL_VEC(INCL_VEC)
  ) mem
  (
    .i_clk                (clk  ),
    .i_reset_n            (reset_n),

    // From EX
    .i_ex_mem_payload     (ex_mem_payload      ),
    .i_ex_mem_vld         (ex_mem_vld          ),

    .i_ex_mem_lqvld_1c    (ex_mem_lqvld_1c     ),
    .i_ex_mem_lqid_1c     (ex_mem_lqid_1c      ),
    .i_ex_mem_lqdata_1c   (ex_mem_lqdata_1c    ),

    .i_ex_mem_lqvld_2c    (ex_mem_lqvld_2c     ),
    .i_ex_mem_lqid_2c     (ex_mem_lqid_2c      ),
    .i_ex_mem_lqdata_2c   (ex_mem_lqdata_2c    ),

    .i_fp_ex_mem_lqvld_1c ('0),
    .i_fp_ex_mem_lqid_1c  ('0),
    .i_fp_ex_mem_lqdata_1c('0),

    .i_fp_ex_mem_lqvld_2c ('0),
    .i_fp_ex_mem_lqid_2c  ('0),
    .i_fp_ex_mem_lqdata_2c('0),

    .i_vex_mem_lqvld_1c   (vex_mem_lqvld_1c),
    .i_vex_mem_lqdata_1c  (vex_mem_lqdata_1c),
    .i_vex_mem_lqexc_1c   (vex_mem_lqexc_1c),
    .i_vex_mem_lqid_1c    (vex_mem_lqid_1c),             
    
    .i_vex_mem_lqvld_2c   (vex_mem_lqvld_2c),
    .i_vex_mem_lqdata_2c  (vex_mem_lqdata_2c),
    .i_vex_mem_lqexc_2c   (vex_mem_lqexc_2c),
    .i_vex_mem_lqid_2c    (vex_mem_lqid_2c),             
    
    .i_vex_mem_lqvld_3c   (vex_mem_lqvld_3c),
    .i_vex_mem_lqdata_3c  (vex_mem_lqdata_3c),
    .i_vex_mem_lqexc_3c   (vex_mem_lqexc_3c),
    .i_vex_mem_lqid_3c    (vex_mem_lqid_3c),             

    // To EX
    .o_mem_ex_rtr         (mem_ex_rtr),

    // To Regfile
    .o_mem_rf_wr          (mem_rf_wr),
    .o_mem_rf_wraddr      (mem_rf_wraddr),
    .o_mem_rf_wrdata      (mem_rf_wrdata),

    //To FP RF
    .o_mem_fp_rf_wr       (mem_fp_rf_wr),
    .o_mem_fp_rf_wraddr   (mem_fp_rf_wraddr),
    .o_mem_fp_rf_wrdata   (mem_fp_rf_wrdata),

    .o_mem_vrf_wr         (mem_vrf_wr),
    .o_mem_vrf_wraddr     (mem_vrf_wraddr),
    .o_mem_vrf_wrdata     (mem_vrf_wrdata),
    .o_mem_vrf_wrexc      (mem_vrf_wrexc),

    .o_vec_store_commit   (vec_store_commit),
    .o_vec_nonstore_commit(vec_nonstore_commit),

    // To ID
    .i_id_mem_lqalloc     (id_mem_lqalloc    ),
    .i_id_mem_lqinfo      (id_mem_lqinfo     ),
    .o_mem_id_lqfull      (mem_fe_lqfull     ),
    .o_mem_id_lqempty     (mem_fe_lqempty     ),
    .o_mem_id_skidbuffull (mem_fe_skidbuffull),
    .o_mem_id_lqnxtid     (mem_id_lqnxtid    ),

    .o_mem_dst_vld        (mem_dst_vld       ),
    .o_mem_dst_lqid       (mem_dst_lqid      ),
    .o_mem_fwd_data       (mem_fwd_data      ),
    .o_mem_lq_op          (mem_lq_op         ),
    .o_mem_lq_commit      (mem_lq_commit     ),

    .o_lq_broadside_info      (lq_broadside_info ),
    .o_lq_broadside_data      (lq_broadside_data ),
    .o_lq_broadside_valid     (lq_broadside_valid),
    .o_lq_broadside_data_valid(lq_broadside_data_valid),

    // To/from memory system
    .i_dmem_brisc_memory_idle('0), 
    .o_data_addr              (o_data_addr       ),
    .o_data_wrdata            (o_wr_data         ),
    .o_data_reqtype           (o_data_reqtype    ),
    .o_data_ordered           (o_data_ordered    ),
    .o_data_byten             (o_data_byten      ), // IMPROVE: rename this signal to reflect its use for loads and stores
    .o_data_req               (o_data_req_prequal),
    .o_data_req_id            (o_data_req_id     ),
    .o_data_128b              (o_data_128b       ),
    .i_data_req_rtr           ('1    ),
    .i_data_vld_0             (load_valid && load_fsm_state == 2   ),
    .i_data_vld_cancel_0      ('0),
    .i_data_resp_id_0         (req_buffer[el_id]),
    .i_data_rddata_0          (load_data[63:0]       ),
    .i_data_vld_1             ('0   ),
    .i_data_vld_cancel_1      ('0),
    .i_data_resp_id_1         ('0),
    .i_data_rddata_1          ('0       ),
    .i_data_vld_2             (i_rd_data_vld_2   ),
    .i_data_vld_cancel_2      ('0),
    .i_data_resp_id_2         (i_rd_data_resp_id_2),
    .i_data_rddata_2          ('0),

    .o_mem_store              (o_mem_store ),
    .o_mem_load               (o_mem_load),
    .o_mem_size               (o_mem_size),
    .o_mem_last               (o_mem_last_raw),
    // Trap
    .i_reset_pc               ('0),
    .o_trap                   (  ),
    .o_lq_empty               (lq_empty)
  );

  logic [LQ_DEPTH     -1:0] lq_last;
  logic [LQ_DEPTH_LOG2-1:0] lq_rd_ptr;

  assign ocelot_instrn_commit_valid       =   mem_rf_wr || mem_fp_rf_wr ||
                                        (vec_nonstore_commit && lq_last[lq_rd_ptr]);
  assign ocelot_instrn_commit_data[VLEN*8-1:64] =  {VLEN*8-64{vec_nonstore_commit}} & mem_vrf_wrdata_nxt[VLEN*8-1:64];
  assign ocelot_instrn_commit_data[      63: 0] =        ({64{vec_nonstore_commit}} & mem_vrf_wrdata_nxt[      63: 0]) |
                                                    ({64{mem_rf_wr          }} & mem_rf_wrdata     [      63: 0]) |
                                                    ({64{mem_fp_rf_wr       }} & mem_fp_rf_wrdata  [      63: 0]);
  assign ocelot_instrn_commit_fflags            =        ({ 5{vec_nonstore_commit}} & mem_vrf_wrexc_nxt [       4: 0]);
  assign ocelot_instrn_commit_mask              =                                     mem_vrf_wrmask_nxt;
  assign o_data_req =  o_data_req_prequal && 
                      !(  o_mem_load   &&
                        ~|o_data_byten   );

  assign o_mem_last = o_mem_last_raw     &&
                      lq_last[o_data_req_id[LQ_DEPTH_LOG2-1:0]];

  always_ff @(posedge clk) begin
    if (!reset_n) begin
        lq_last          <= '0;
        lq_rd_ptr        <= '0;
        mem_id_lqnxtid_r <= '0;
    end else begin
        if (mem_lq_commit) begin
          lq_rd_ptr <= lq_rd_ptr + 1;
        end

        if (id_mem_lqalloc) begin
          lq_last[mem_id_lqnxtid] <= id_mem_lq_done;
          mem_id_lqnxtid_r        <= mem_id_lqnxtid;
        end else
        if (id_mem_lq_done) begin
          lq_last[mem_id_lqnxtid_r] <= 1'b1;
        end
    end
  end


  logic [2:0] lmul_cnt;

  always_ff @(posedge clk) begin
    if (!reset_n) begin
        mem_vrf_wrdata_reg <= '0;
        mem_vrf_wrmask_reg <= '0;
        mem_vrf_wrexc_reg  <= '0;
    end else begin
        if (ocelot_instrn_commit_valid) begin
          mem_vrf_wrdata_reg <= '0;
          mem_vrf_wrmask_reg <= '0;
          mem_vrf_wrexc_reg  <= '0;
        end else
        if (mem_vrf_wr) begin
          mem_vrf_wrdata_reg <= mem_vrf_wrdata_nxt;
          mem_vrf_wrmask_reg <= mem_vrf_wrmask_nxt;
          mem_vrf_wrexc_reg  <= mem_vrf_wrexc_nxt;
        end
    end
  end

  always_comb begin
    mem_vrf_wrdata_nxt = mem_vrf_wrdata_reg;
    mem_vrf_wrmask_nxt = mem_vrf_wrmask_reg;
    mem_vrf_wrexc_nxt  = mem_vrf_wrexc_reg;

    mem_vrf_wrdata_nxt[VLEN*lmul_cnt +: VLEN] = mem_vrf_wrdata;
    mem_vrf_wrmask_nxt[     lmul_cnt        ] = |vcsr[$clog2(VLEN+1)-1+14:14];
    mem_vrf_wrexc_nxt                        |= mem_vrf_wrexc;
  end

  always_ff @(posedge clk) begin
    if (!reset_n) begin
        lmul_cnt <= '0;
    end else begin
        if (ocelot_instrn_commit_valid) begin
          lmul_cnt <= '0;
        end else
        if (mem_vrf_wr) begin
          lmul_cnt <= lmul_cnt + 1;
        end
    end
  end

  always_ff @(posedge clk) begin
    if (!reset_n) begin
        i_rd_data_vld_2 <= '0;
        i_rd_data_resp_id_2 <= '0;
    end else begin
        i_rd_data_vld_2 <=   o_data_req_prequal &&
                            '1     &&
                          (  o_mem_load   &&
                            ~|o_data_byten   );
        i_rd_data_resp_id_2 <= o_data_req_id;
    end
  end

  assign enough_data = store_buffer_valid[store_buffer_rptr] && !store_buffer_sent[store_buffer_rptr] &&
                       store_buffer_valid[store_buffer_rptr+1] && !store_buffer_sent[store_buffer_rptr+1];
  always_comb begin
    store_fsm_next_state = 0;
    case (store_fsm_state)
      0: begin
        if(vecldst_autogen_store && ocelot_read_req) begin
          if(id_mem_lq_done)
            store_fsm_next_state = 2;
          else
            store_fsm_next_state = 1;
        end
      end

      1: begin
        if(id_mem_lq_done)
          store_fsm_next_state = 2;
        else
          store_fsm_next_state = 1;
      end

      2: begin
        if(memop_sync_end)
          store_fsm_next_state = 3;
        else
          store_fsm_next_state = 2;
      end

      3: begin
        if(lq_empty)
          store_fsm_next_state = 0;
        else
          store_fsm_next_state = 3;
      end
    endcase
  end

  always_ff@(posedge clk) begin
    if(!reset_n) begin
      store_buffer_wptr <= 0;
      store_fsm_state <= 0;
      store_buffer_full <= 0;
      store_credits <= STORE_CREDITS;
    end
    else begin
      store_fsm_state <= store_fsm_next_state;

      // Reset the store buffer when idle
      if(store_fsm_state == 0 && !vecldst_autogen_store) begin
        for(int i=0; i<8; i=i+1)
          store_buffer[i] <= 0;
        store_buffer_full <= 0;
        store_buffer_valid <= 0;
        store_buffer_wptr <= 0;
      end
      else if(store_fsm_state == 1 || (store_fsm_state == 0 && vecldst_autogen_store && ocelot_read_req)) begin
        if(id_ex_units_rts) begin
          store_buffer[store_buffer_wptr] <= vs3_rddata;
          store_buffer_valid[store_buffer_wptr] <= 1;
          store_buffer_wptr <= store_buffer_wptr + 1;
          if(store_buffer_wptr == 7)
            store_buffer_full <= 1;
        end
      end
    end
  end

  assign store_memsync_start = store_fsm_state == 0 && vecldst_autogen_store && ocelot_read_req;
  always_ff@(posedge clk) begin
    if(!reset_n)
      memop_sync_start <= 0;
    else
      memop_sync_start <= store_memsync_start | load_memsync_start;
  end

  always_ff@(posedge clk) begin
    if(!reset_n) begin
      store_valid <= 0;
      store_data <= 0;
      store_commit <= 0;
      store_buffer_rptr <= 0;
      store_buffer_sent <= 0;
    end
    else begin
      if((store_fsm_state == 0 || store_fsm_next_state == 0) && !vecldst_autogen_store) begin
        store_buffer_rptr <= 0;
        store_buffer_sent <= 0;
      end
      // Bypass the store buffer because we only need to send 1 register
      else if((store_fsm_state == 1 || store_fsm_state == 0) && id_ex_units_rts && vecldst_autogen_store && ocelot_read_req && id_mem_lq_done && store_buffer_wptr == 0) begin
        store_valid <= 1;
        store_data[255:0] <= vs3_rddata;
      end
      else if((store_fsm_state == 1 || store_fsm_state == 2) && enough_data && store_credits > 0) begin
        store_valid <= 1;
        // little endian
        store_data[255:0] <= store_buffer[store_buffer_rptr];
        store_data[511:256] <= store_buffer[store_buffer_rptr+1];
        store_buffer_sent[store_buffer_rptr] <= 1;
        store_buffer_sent[store_buffer_rptr+1] <= 1;
        store_buffer_rptr <= store_buffer_rptr + 2;
      end
      else
        store_valid <= 0;

      if(store_fsm_state == 3 && lq_empty)
        store_commit <= 1;
      else
        store_commit <= 0;
    end
  end

  // This queue should never overflow, so I'm not going to add phase bits
  // to check if it's full or not.
  localparam sbid_queue_depth = 8;
  logic [sbid_queue_depth-1:0][4:0] sbid_queue;
  logic [$clog2(sbid_queue_depth)-1:0] sbid_queue_wptr;
  logic [$clog2(sbid_queue_depth)-1:0] sbid_queue_rptr;

  always_ff@(posedge clk) begin
    if(!reset_n) begin
      for(int i=0; i<sbid_queue_depth; i=i+1)
        sbid_queue[i] <= 0;
      sbid_queue_wptr <= 0;
      sbid_queue_rptr <= 0;
    end
    else begin
      if(ocelot_read_req && read_valid) begin
        sbid_queue[sbid_queue_wptr] <= read_issue_sb_id;
        sbid_queue_wptr <= sbid_queue_wptr + 1;
      end
      if((ocelot_instrn_commit_valid && load_fsm_state != 2'd2) || store_commit || load_commit) begin
        sbid_queue_rptr <= sbid_queue_rptr + 1;
      end
    end
  end

  assign issue_credit = 0;

  tt_fifo #(
    .DEPTH(16)
  ) fifo0
  (
    .clk(clk),
    .reset_n(reset_n),

    .issue_inst(issue_inst),
    .issue_sb_id(issue_sb_id),
    .issue_scalar_opnd(issue_scalar_opnd),
    .issue_vcsr(issue_vcsr),
    .issue_vcsr_lmulb2(issue_vcsr_lmulb2),
    .issue_valid(issue_valid),

    .dispatch_sb_id(dispatch_sb_id),
    .dispatch_next_senior(dispatch_next_senior),
    .dispatch_kill(dispatch_kill),

    .read_req(ocelot_read_req),
    .read_valid(read_valid),
    .read_issue_inst(read_issue_inst),
    .read_issue_sb_id(read_issue_sb_id),
    .read_issue_scalar_opnd(read_issue_scalar_opnd),
    .read_issue_vcsr(read_issue_vcsr),
    .read_issue_vcsr_lmulb2(read_issue_vcsr_lmulb2)
  );

  assign vcsr        = ocelot_read_req && read_valid ? read_issue_vcsr : vcsr_reg;
  assign vcsr_lmulb2 = ocelot_read_req && read_valid ? read_issue_vcsr_lmulb2 : vcsr_lmulb2_reg;

  always_ff@(posedge clk) begin
    if(!reset_n)
      {vcsr_reg, vcsr_lmulb2_reg} <= 0;
    else if(read_valid && ocelot_read_req) begin
      vcsr_reg <= read_issue_vcsr;
      vcsr_lmulb2_reg <= read_issue_vcsr_lmulb2;
    end
  end

  assign v_reg = load_seq_id[4:0];
  assign el_id = load_seq_id[15:5];
  assign el_off = load_seq_id[21:16];
  assign el_count = load_seq_id[28:22];
  assign sb_id = load_seq_id[33:29];

  always @(posedge clk) begin
    if(!reset_n)
      {eew,load_stride,eew_log2} <= 0;
    else if(read_valid && ocelot_read_req) begin
      eew <= read_issue_inst[14:12] == 3'b000 ? 2'd0 : // 8-bit EEW
             read_issue_inst[14:12] == 3'b101 ? 2'd1 : // 16-bit EEW
             read_issue_inst[14:12] == 3'b110 ? 2'd2 : 2'd3; // 32-bit, 64-bit EEW
      eew_log2 <= read_issue_inst[14:12] == 3'b000 ? 3'd3 : // 8-bit EEW
                  read_issue_inst[14:12] == 3'b101 ? 3'd4 : // 16-bit EEW
                  read_issue_inst[14:12] == 3'b110 ? 3'd5 : 3'd6; // 32-bit, 64-bit EEW
      load_stride <= read_issue_scalar_opnd;
    end
  end

  integer i,j;
  always_comb begin
    packed_load_data = load_data;
    case(eew)
      2'd0: begin
        case($signed(load_stride))
          64'd1: begin 
            packed_load_data = load_data;
            load_stride_in_eew_log2 = 0;
          end
          -64'd1: begin
            for(i=0, j=511; i<512; i=i+8, j=j-8)
              packed_load_data[i+:8] = load_data[j-:8];
            load_stride_in_eew_log2 = 0;
          end
          64'd2: begin
            for(i=0, j=0; i<256; i=i+8, j=j+16)
              packed_load_data[i+:8] = el_off[0] ? load_data[j+8+:8] : load_data[j+:8];
            load_stride_in_eew_log2 = 1;
          end
          -64'd2: begin
            for(i=0, j=511; i<256; i=i+8, j=j-16)
              packed_load_data[i+:8] = el_off[0] ? load_data[j-8-:8] : load_data[j-:8];
            load_stride_in_eew_log2 = 1;
          end
          64'd4: begin
            for(i=0, j=0; i<128; i=i+8, j=j+32)
              packed_load_data[i+:8] = el_off[1:0] == 2'b00 ? load_data[j+:8] :
                                         el_off[1:0] == 2'b01 ? load_data[j+8+:8] :
                                         el_off[1:0] == 2'b10 ? load_data[j+16+:8] : load_data[j+23+:8];
            load_stride_in_eew_log2 = 2;
          end
          -64'd4: begin
            for(i=0, j=511; i<128; i=i+8, j=j-32)
              packed_load_data[i+:8] = el_off[1:0] == 2'b00 ? load_data[j-:8] :
                                         el_off[1:0] == 2'b01 ? load_data[j-8-:8] :
                                         el_off[1:0] == 2'b10 ? load_data[j-16-:8] : load_data[j-23-:8];
            load_stride_in_eew_log2 = 2;
          end
        endcase
      end
      2'd1: begin
      case($signed(load_stride))
        64'd2: begin 
          packed_load_data = load_data;
          load_stride_in_eew_log2 = 0;
        end
        -64'd2: begin
          for(i=0, j=511; i<512; i=i+16, j=j-16)
            packed_load_data[i+:16] = load_data[j-:16];
          load_stride_in_eew_log2 = 0;
        end
        64'd4: begin
          for(i=0, j=0; i<256; i=i+16, j=j+32)
            packed_load_data[i+:16] = el_off[0] ? load_data[j+16+:16] : load_data[j+:16];
          load_stride_in_eew_log2 = 1;
        end
        -64'd4: begin
          for(i=0, j=511; i<256; i=i+16, j=j-32)
            packed_load_data[i+:16] = el_off[0] ? load_data[j-16-:16] : load_data[j-:16];
          load_stride_in_eew_log2 = 1;
        end
        64'd8: begin
          for(i=0, j=0; i<128; i=i+16, j=j+64)
            packed_load_data[i+:16] = el_off[1:0] == 2'b00 ? load_data[j+:16] :
                                      el_off[1:0] == 2'b01 ? load_data[j+16+:16] :
                                      el_off[1:0] == 2'b10 ? load_data[j+32+:16] : load_data[j+48+:16];
          load_stride_in_eew_log2 = 2;
        end
        -64'd8: begin
          for(i=0, j=511; i<128; i=i+16, j=j-64)
            packed_load_data[i+:16] = el_off[1:0] == 2'b00 ? load_data[j-:16] :
                                      el_off[1:0] == 2'b01 ? load_data[j-16-:16] :
                                      el_off[1:0] == 2'b10 ? load_data[j-32-:16] : load_data[j-48-:16];
          load_stride_in_eew_log2 = 2;
        end
      endcase
      end
      2'd2: begin
      case($signed(load_stride))
        64'd4: begin 
          packed_load_data = load_data;
          load_stride_in_eew_log2 = 0;
        end
        -64'd4: begin
          for(i=0, j=511; i<512; i=i+32, j=j-32)
            packed_load_data[i+:32] = load_data[j-:32];
          load_stride_in_eew_log2 = 0;
        end
        64'd8: begin
          for(i=0, j=0; i<256; i=i+32, j=j+64)
            packed_load_data[i+:32] = el_off[0] ? load_data[j+63-:32] : load_data[j+31-:32];
          load_stride_in_eew_log2 = 1;
        end
        -64'd8: begin
          for(i=0, j=511; i<256; i=i+32, j=j-64)
            packed_load_data[i+:32] = el_off[0] ? load_data[j-32-:32] : load_data[j-:32];
          load_stride_in_eew_log2 = 1;
        end
        64'd16: begin
          for(i=0, j=0; i<128; i=i+32, j=j+128)
            packed_load_data[i+:32] = el_off[1:0] == 2'b00 ? load_data[j+31-:32] :
                                      el_off[1:0] == 2'b01 ? load_data[j+63-:32] :
                                      el_off[1:0] == 2'b10 ? load_data[j+95-:32] : load_data[j+127-:32];
          load_stride_in_eew_log2 = 2;
        end
        -64'd16: begin
          for(i=0, j=511; i<128; i=i+32, j=j-128)
            packed_load_data[i+:32] = el_off[1:0] == 2'b00 ? load_data[j-:32] :
                                      el_off[1:0] == 2'b01 ? load_data[j-32-:32] :
                                      el_off[1:0] == 2'b10 ? load_data[j-64-:32] : load_data[j-96-:32];
          load_stride_in_eew_log2 = 2;
        end
      endcase
      end
      2'd3: begin
      case($signed(load_stride))
        64'd8: begin
          packed_load_data = load_data;
          load_stride_in_eew_log2 = 0;
        end
        -64'd8: begin
          for(i=0, j=511; i<512; i=i+64, j=j-64)
            packed_load_data[i+:64] = load_data[j-:64];
          load_stride_in_eew_log2 = 0;
        end
        64'd16: begin
          for(i=0, j=0; i<256; i=i+64, j=j+128)
            packed_load_data[i+:64] = el_off[0] ? load_data[j+127-:64] : load_data[j+63-:64];
          load_stride_in_eew_log2 = 1;
        end
        -64'd16: begin
          for(i=0, j=511; i<256; i=i+64, j=j-128)
            packed_load_data[i+:64] = el_off[0] ? load_data[j-64-:64] : load_data[j-:64];
          load_stride_in_eew_log2 = 1;
        end
        64'd32: begin
          for(i=0, j=0; i<128; i=i+64, j=j+256)
            packed_load_data[i+:64] = el_off[1:0] == 2'b00 ? load_data[j+63-:64] :
                                      el_off[1:0] == 2'b01 ? load_data[j+127-:64] :
                                      el_off[1:0] == 2'b10 ? load_data[j+191-:64] : load_data[j+255-:64];
          load_stride_in_eew_log2 = 2;
        end
        -64'd32: begin
          for(i=0, j=511; i<128; i=i+64, j=j-256)
            packed_load_data[i+:64] = el_off[1:0] == 2'b00 ? load_data[j-:64] :
                                      el_off[1:0] == 2'b01 ? load_data[j-64-:64] :
                                      el_off[1:0] == 2'b10 ? load_data[j-128-:64] : load_data[j-192-:64];
          load_stride_in_eew_log2 = 2;
        end
      endcase
      end
    endcase
  end

  always_comb begin
    packed_offset = el_off >> load_stride_in_eew_log2;
    offset_diff = (el_id - packed_offset) << eew_log2;
    shamt = offset_diff[10] ? offset_diff + VLEN : offset_diff;
    // Circular rotate left by shamt
    // shifted_load_data = packed_load_data << shamt | (packed_load_data >> (512-shamt));
    shifted_load_data = packed_load_data << (el_id << eew_log2);
    el_id_lower_bound = el_id << eew_log2;
    el_id_upper_bound = (el_id + el_count) << eew_log2;
  end

  integer k;
  always @(posedge clk) begin
    if(!reset_n)
      for(k=0; k<8; k=k+1)
        load_buffer[k] <= 0;
    else begin
      for(k=0; k<VLEN; k=k+1)
        load_buffer[v_reg[2:0]][k] <= (el_id_lower_bound <= k && k < el_id_upper_bound) ? shifted_load_data[k] : load_buffer[v_reg[2:0]][k];
    end
  end

  always_comb begin
    load_fsm_next_state = 2'd0;
    case(load_fsm_state)
      2'd0: begin
        if(vecldst_autogen_load && ocelot_read_req)
          load_fsm_next_state = 2'd1;
        else
          load_fsm_next_state = 2'd0;
      end
      2'd1: begin
        if(!o_data_req && req_buffer_wptr != 0)
          load_fsm_next_state = 2'd2;
        else
          load_fsm_next_state = 2'd1;
      end
      2'd2: begin
        if(memop_sync_end)
          load_fsm_next_state = 2'd3;
        else
          load_fsm_next_state = 2'd2;
      end
      2'd3: begin
        if(lq_empty)
          load_fsm_next_state = 2'd0;
        else
          load_fsm_next_state = 2'd3;
      end
    endcase
  end
  assign load_memsync_start = load_fsm_state == 2'd1 && load_fsm_next_state == 2'd2;
  assign load_commit = load_fsm_state == 2'd3 && lq_empty;

  assign ovi_stall = store_fsm_state != 0 || load_fsm_state != 0;

  always_ff@(posedge clk) begin
    if(!reset_n)
      load_fsm_state <= 0;
    else
      load_fsm_state <= load_fsm_next_state;
  end

  integer r;
  always @(posedge clk) begin
    if(!reset_n) begin
      req_buffer_wptr <= 0;
      for(r=0; r<VLEN; r=r+1)
        req_buffer[r] <= 0;
    end
    else begin
      if(load_fsm_state == 0) begin
        req_buffer_wptr <= 0;
        for(r=0; r<VLEN; r=r+1)
          req_buffer[r] <= 0;
      end
      else if(load_fsm_state == 1 && o_data_req) begin
        req_buffer[req_buffer_wptr] <= o_data_req_id;
        req_buffer_wptr <= req_buffer_wptr + 1;
      end
    end
  end


  // Just pass the parameters down...
  // vfp_pipeline #(
  //   .LOCAL_MEM_BYTE_ADDR_WIDTH(LOCAL_MEM_BYTE_ADDR_WIDTH),
  //   .INCL_VEC(INCL_VEC),
  //   .VLEN(VLEN),
  //   .ADDRWIDTH(ADDRWIDTH),
  //   .LD_DATA_WIDTH_BITS(LD_DATA_WIDTH_BITS),
  //   .ST_DATA_WIDTH_BITS(ST_DATA_WIDTH_BITS),
  //   .LQ_DEPTH(LQ_DEPTH),
  //   .LQ_DEPTH_LOG2(LQ_DEPTH_LOG2),
  //   .DATA_REQ_ID_WIDTH(DATA_REQ_ID_WIDTH),
  //   .INCL_FP(INCL_FP)
  // ) ocelot
  // (
  //   .i_clk(clk),
  //   .i_reset(!reset_n),
  //   .i_csr_vl(vcsr[$clog2(VLEN+1)-1+14:14]),
  //   .i_csr_vsew(vcsr[38:36]),
  //   .i_csr_vlmul({vcsr_lmulb2,vcsr[35:34]}),
  //   .i_csr_vxrm(vcsr[30:29]),
  //   .i_csr_frm(vcsr[33:31]),

  //   // IF Interface
  //   .i_if_instrn_rts(read_valid),
  //   .o_id_instrn_rtr(ocelot_read_req),
  //   .i_if_instrn(read_issue_inst),
  //   .i_if_pc(0),
  //   .i_rf_vex_p0(read_issue_scalar_opnd),
  //   .i_rf_vex_p1(read_issue_scalar_opnd),
  //   .i_fprf_vex_p0(read_issue_scalar_opnd),

  //   // Commit Interface
  //   .o_instrn_commit_valid(ocelot_instrn_commit_valid),
  //   .o_instrn_commit_data(ocelot_instrn_commit_data),
  //   .o_instrn_commit_mask(ocelot_instrn_commit_mask),
  //   .o_instrn_commit_fflags(ocelot_instrn_commit_fflags),

  //   .o_sat_csr(ocelot_sat_csr),

  //   // Memory Interface
  //   .o_data_req(o_data_req),
  //   .o_data_addr(o_data_addr),
  //   .o_data_byten(o_data_byten),
  //   .o_wr_data(o_wr_data),
  //   .o_data_req_id(o_data_req_id),
  //   .o_mem_load(o_mem_load),
  //   .o_mem_size(o_mem_size),
  //   .o_mem_last(o_mem_last),
  //   .i_data_req_rtr('1),
  //   .i_rd_data_vld_0(load_valid && load_fsm_state == 2),
  //   .i_rd_data_resp_id_0(req_buffer[el_id]),
  //   .i_rd_data_0(load_data[63:0]),
  //   .i_rd_data_vld_1('0),
  //   .i_rd_data_resp_id_1('0),
  //   .i_rd_data_1('0),

  //   .o_vecldst_autogen_store(vecldst_autogen_store),
  //   .o_vecldst_autogen_load(vecldst_autogen_load),
  //   .o_id_mem_lq_done(id_mem_lq_done),
  //   .o_id_ex_units_rts(id_ex_units_rts),
  //   .o_vs3_rddata(vs3_rddata),
  //   .o_lq_empty(lq_empty),

  //   .i_ovi_stall(ovi_stall)
  // );

  always @(posedge clk) begin
    if(!reset_n) begin
      completed_valid <= 0;
      completed_sb_id <= 0;
      completed_fflags <= 0;
      completed_dest_reg <= 0;
      completed_vxsat <= 0;
      completed_vstart <= 0;
      completed_illegal <= 0;
    end
    else begin
      completed_valid <= (ocelot_instrn_commit_valid && load_fsm_state != 2'd2) || store_commit || load_commit;
      completed_sb_id <= sbid_queue[sbid_queue_rptr];
      completed_fflags <= ocelot_instrn_commit_fflags;
      completed_dest_reg <= ocelot_instrn_commit_data[63:0];
      completed_vxsat <= 0;
      completed_vstart <= 0;
      completed_illegal <= 0;
    end
  end

  assign debug_wb_vec_valid = ocelot_instrn_commit_valid;
  assign debug_wb_vec_wdata = ocelot_instrn_commit_data;
  assign debug_wb_vec_wmask = ocelot_instrn_commit_mask;

endmodule
