// See LICENSE.TT for license details.

// Allow multiple modules in autogen file
//spyglass disable_block OneModule-ML
// Cases can sometimes overlap for specific values, but that is fine
//spyglass disable_block W398

module autogen_Instruction (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [0:0] vm,
input [2:0] sew,
input [2:0] lmul,
input [1:0] mop,
input [4:0] SrcB,
input [2:0] nf,
output reg [127:0] Instruction
);
//spyglass disable_block STARC05-2.10.3.2b_sa
//spyglass disable_block STARC05-2.10.3.2b_sb
//spyglass disable_block W164c

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0], vm[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0], nf[2], nf[1], nf[0]})
	    34'b1110011???????001?????????????????  :  Instruction = "CSRRW";
	    34'b1110011???????010?????????????????  :  Instruction = "CSRRS";
	    34'b1110011???????011?????????????????  :  Instruction = "CSRRC";
	    34'b1110011???????101?????????????????  :  Instruction = "CSRRWI";
	    34'b1110011???????110?????????????????  :  Instruction = "CSRRSI";
	    34'b1110011???????111?????????????????  :  Instruction = "CSRRCI";
	    34'b0110111???????????????????????????  :  Instruction = "LUI";
	    34'b0010111???????????????????????????  :  Instruction = "AUIPC";
	    34'b1101111???????????????????????????  :  Instruction = "JAL";
	    34'b1100111???????000?????????????????  :  Instruction = "JALR";
	    34'b1100011???????000?????????????????  :  Instruction = "BEQ";
	    34'b1100011???????001?????????????????  :  Instruction = "BNE";
	    34'b1100011???????100?????????????????  :  Instruction = "BLT";
	    34'b1100011???????101?????????????????  :  Instruction = "BGE";
	    34'b1100011???????110?????????????????  :  Instruction = "BLTU";
	    34'b1100011???????111?????????????????  :  Instruction = "BGEU";
	    34'b0000011???????000?????????????????  :  Instruction = "LB";
	    34'b0000011???????001?????????????????  :  Instruction = "LH";
	    34'b0000011???????010?????????????????  :  Instruction = "LW";
	    34'b0000011???????100?????????????????  :  Instruction = "LBU";
	    34'b0000011???????101?????????????????  :  Instruction = "LHU";
	    34'b0100011???????000?????????????????  :  Instruction = "SB";
	    34'b0100011???????001?????????????????  :  Instruction = "SH";
	    34'b0100011???????010?????????????????  :  Instruction = "SW";
	    34'b0010011???????000?????????????????  :  Instruction = "ADDI";
	    34'b0010011???????010?????????????????  :  Instruction = "SLTI";
	    34'b0010011???????011?????????????????  :  Instruction = "SLTIU";
	    34'b0010011???????100?????????????????  :  Instruction = "XORI";
	    34'b0010011???????110?????????????????  :  Instruction = "ORI";
	    34'b0010011???????111?????????????????  :  Instruction = "ANDI";
	    34'b00100110000000001?????????????????  :  Instruction = "SLLI";
	    34'b00100110000000101?????????????????  :  Instruction = "SRLI";
	    34'b00100110100000101?????????????????  :  Instruction = "SRAI";
	    34'b01100110000000000?????????????????  :  Instruction = "ADD";
	    34'b01100110100000000?????????????????  :  Instruction = "SUB";
	    34'b01100110000000001?????????????????  :  Instruction = "SLL";
	    34'b01100110000000010?????????????????  :  Instruction = "SLT";
	    34'b01100110000000011?????????????????  :  Instruction = "SLTU";
	    34'b01100110000000100?????????????????  :  Instruction = "XOR";
	    34'b01100110000000101?????????????????  :  Instruction = "SRL";
	    34'b01100110100000101?????????????????  :  Instruction = "SRA";
	    34'b01100110000000110?????????????????  :  Instruction = "OR";
	    34'b01100110000000111?????????????????  :  Instruction = "AND";
	    34'b0001111???????000?????????????????  :  Instruction = "FENCE";
	    34'b1110011???????000?????????????????  :  Instruction = "ECALL";
	    34'b00000000000000000?????????????????  :  Instruction = "ILLEGAL";
	    34'b01100110000001000?????????????????  :  Instruction = "MUL";
	    34'b01100110000001001?????????????????  :  Instruction = "MULH";
	    34'b01100110000001010?????????????????  :  Instruction = "MULHSU";
	    34'b01100110000001011?????????????????  :  Instruction = "MULHU";
	    34'b01100110000001100?????????????????  :  Instruction = "DIV";
	    34'b01100110000001101?????????????????  :  Instruction = "DIVU";
	    34'b01100110000001110?????????????????  :  Instruction = "REM";
	    34'b01100110000001111?????????????????  :  Instruction = "REMU";
	    34'b010111100001??010?????????????????  :  Instruction = "AMOSWAP";
	    34'b0101111000????010?????????????????  :  Instruction = "AMOADD";
	    34'b0101111001????010?????????????????  :  Instruction = "AMOXOR";
	    34'b0101111010????010?????????????????  :  Instruction = "AMOAND";
	    34'b0101111011????010?????????????????  :  Instruction = "AMOOR";
	    34'b0101111100????010?????????????????  :  Instruction = "AMOMIN";
	    34'b0101111101????010?????????????????  :  Instruction = "AMOMAX";
	    34'b0101111110????010?????????????????  :  Instruction = "AMOMINU";
	    34'b0101111111????010?????????????????  :  Instruction = "AMOMAXU";
	    34'b00100110110000001?????????????????  :  Instruction = "CLZ";
	    34'b01100110000101100?????????????????  :  Instruction = "MIN";
	    34'b01100110000101101?????????????????  :  Instruction = "MINU";
	    34'b01100110000101110?????????????????  :  Instruction = "MAX";
	    34'b01100110000101111?????????????????  :  Instruction = "MAXU";
	    34'b01100110000100100?????????????????  :  Instruction = "PACK";
	    34'b01100110100000111?????????????????  :  Instruction = "ANDN";
	    34'b01100110100000110?????????????????  :  Instruction = "ORN";
	    34'b01100110100000100?????????????????  :  Instruction = "XNOR";
	    34'b01100110110000001?????????????????  :  Instruction = "ROL";
	    34'b01100110110000101?????????????????  :  Instruction = "ROR";
	    34'b001001101100??101?????????????????  :  Instruction = "RORI";
	    34'b001001101101??101?????????????????  :  Instruction = "GREVI";
	    34'b001001100101??101?????????????????  :  Instruction = "GORCI";
	    34'b01100110010000010?????????????????  :  Instruction = "SH1ADD";
	    34'b01100110010000100?????????????????  :  Instruction = "SH2ADD";
	    34'b01100110010000110?????????????????  :  Instruction = "SH3ADD";
	    34'b0000111???????010?????????????????  :  Instruction = "FLW";
	    34'b0100111???????010?????????????????  :  Instruction = "FSW";
	    34'b10100110000000????????????????????  :  Instruction = "FADD.S";
	    34'b10100110000100????????????????????  :  Instruction = "FSUB.S";
	    34'b10100110001000????????????????????  :  Instruction = "FMUL.S";
	    34'b10100110010100000?????????????????  :  Instruction = "FMIN.S";
	    34'b10100110010100001?????????????????  :  Instruction = "FMAX.S";
	    34'b1000011?????00????????????????????  :  Instruction = "FMADD.S";
	    34'b1000111?????00????????????????????  :  Instruction = "FMSUB.S";
	    34'b1001111?????00????????????????????  :  Instruction = "FNMADD.S";
	    34'b1001011?????00????????????????????  :  Instruction = "FNMSUB.S";
	    34'b10100111100000????????????????????  :  Instruction = "FCVT.W.S";
	    34'b10100111101000????????????????????  :  Instruction = "FCVT.S.W";
	    34'b10100110010000000?????????????????  :  Instruction = "FSGNJ.S";
	    34'b10100110010000001?????????????????  :  Instruction = "FSGNJN.S";
	    34'b10100110010000010?????????????????  :  Instruction = "FSGNJX.S";
	    34'b10100111110000000?????????????????  :  Instruction = "FMV.X.W";
	    34'b10100111111000000?????????????????  :  Instruction = "FMV.W.X";
	    34'b10100111010000010?????????????????  :  Instruction = "FEQ.S";
	    34'b10100111010000001?????????????????  :  Instruction = "FLT.S";
	    34'b10100111010000000?????????????????  :  Instruction = "FLE.S";
	    34'b10100111110000001?????????????????  :  Instruction = "FCLASS.S";
	    34'b0000111???????001?????????????????  :  Instruction = "FLH";
	    34'b0100111???????001?????????????????  :  Instruction = "FSH";
	    34'b10100110000010????????????????????  :  Instruction = "FADD.H";
	    34'b10100110000110????????????????????  :  Instruction = "FSUB.H";
	    34'b10100110001010????????????????????  :  Instruction = "FMUL.H";
	    34'b10100110010110000?????????????????  :  Instruction = "FMIN.H";
	    34'b10100110010110001?????????????????  :  Instruction = "FMAX.H";
	    34'b1000011?????10????????????????????  :  Instruction = "FMADD.H";
	    34'b1000111?????10????????????????????  :  Instruction = "FMSUB.H";
	    34'b1001111?????10????????????????????  :  Instruction = "FNMADD.H";
	    34'b1001011?????10????????????????????  :  Instruction = "FNMSUB.H";
	    34'b10100111100010????????????????????  :  Instruction = "FCVT.W.H";
	    34'b10100111101010????????????????????  :  Instruction = "FCVT.H.W";
	    34'b10100110100010????????????????????  :  Instruction = "FCVT.H.S";
	    34'b10100110100000????????????????????  :  Instruction = "FCVT.S.H";
	    34'b10100110010010000?????????????????  :  Instruction = "FSGNJ.H";
	    34'b10100110010010001?????????????????  :  Instruction = "FSGNJN.H";
	    34'b10100110010010010?????????????????  :  Instruction = "FSGNJX.H";
	    34'b10100111110010000?????????????????  :  Instruction = "FMV.X.H";
	    34'b10100111111010000?????????????????  :  Instruction = "FMV.H.X";
	    34'b10100111010010010?????????????????  :  Instruction = "FEQ.H";
	    34'b10100111010010001?????????????????  :  Instruction = "FLT.H";
	    34'b10100111010010000?????????????????  :  Instruction = "FLE.H";
	    34'b10100111110010001?????????????????  :  Instruction = "FCLASS.H";
	    34'b10101110??????111?????????????????  :  Instruction = "VSETVLI";
	    34'b101011111?????111?????????????????  :  Instruction = "VSETIVLI";
	    34'b1010111100000?111?????????????????  :  Instruction = "VSETVL";
	    34'b1010111000000?000?????????????????  :  Instruction = "VADD.vv";
	    34'b1010111000000?100?????????????????  :  Instruction = "VADD.vx";
	    34'b1010111000000?011?????????????????  :  Instruction = "VADD.vi";
	    34'b1010111000010?000?????????????????  :  Instruction = "VSUB.vv";
	    34'b1010111000010?100?????????????????  :  Instruction = "VSUB.vx";
	    34'b1010111000011?100?????????????????  :  Instruction = "VRSUB.vx";
	    34'b1010111000011?011?????????????????  :  Instruction = "VRSUB.vi";
	    34'b1010111110000?010?????????????????  :  Instruction = "VWADDU.vv";
	    34'b1010111110000?110?????????????????  :  Instruction = "VWADDU.vx";
	    34'b1010111110010?010?????????????????  :  Instruction = "VWSUBU.vv";
	    34'b1010111110010?110?????????????????  :  Instruction = "VWSUBU.vx";
	    34'b1010111110001?010?????????????????  :  Instruction = "VWADD.vv";
	    34'b1010111110001?110?????????????????  :  Instruction = "VWADD.vx";
	    34'b1010111110011?010?????????????????  :  Instruction = "VWSUB.vv";
	    34'b1010111110011?110?????????????????  :  Instruction = "VWSUB.vx";
	    34'b1010111110100?010?????????????????  :  Instruction = "VWADDU.wv";
	    34'b1010111110100?110?????????????????  :  Instruction = "VWADDU.wx";
	    34'b1010111110110?010?????????????????  :  Instruction = "VWSUBU.wv";
	    34'b1010111110110?110?????????????????  :  Instruction = "VWSUBU.wx";
	    34'b1010111110101?010?????????????????  :  Instruction = "VWADD.wv";
	    34'b1010111110101?110?????????????????  :  Instruction = "VWADD.wx";
	    34'b1010111110111?010?????????????????  :  Instruction = "VWSUB.wv";
	    34'b1010111110111?110?????????????????  :  Instruction = "VWSUB.wx";
	    34'b1010111010000?0000????????????????  :  Instruction = "VADC.vvm";
	    34'b1010111010000?1000????????????????  :  Instruction = "VADC.vxm";
	    34'b1010111010000?0110????????????????  :  Instruction = "VADC.vim";
	    34'b1010111010001?0000????????????????  :  Instruction = "VMADC.vvm";
	    34'b1010111010001?1000????????????????  :  Instruction = "VMADC.vxm";
	    34'b1010111010001?0110????????????????  :  Instruction = "VMADC.vim";
	    34'b1010111010001?000?????????????????  :  Instruction = "VMADC.vv";
	    34'b1010111010001?100?????????????????  :  Instruction = "VMADC.vx";
	    34'b1010111010001?011?????????????????  :  Instruction = "VMADC.vi";
	    34'b1010111010010?0000????????????????  :  Instruction = "VSBC.vvm";
	    34'b1010111010010?1000????????????????  :  Instruction = "VSBC.vxm";
	    34'b1010111010011?0000????????????????  :  Instruction = "VMSBC.vvm";
	    34'b1010111010011?1000????????????????  :  Instruction = "VMSBC.vxm";
	    34'b1010111010011?0001????????????????  :  Instruction = "VMSBC.vv";
	    34'b1010111010011?1001????????????????  :  Instruction = "VMSBC.vx";
	    34'b1010111001001?000?????????????????  :  Instruction = "VAND.vv";
	    34'b1010111001001?100?????????????????  :  Instruction = "VAND.vx";
	    34'b1010111001001?011?????????????????  :  Instruction = "VAND.vi";
	    34'b1010111001010?000?????????????????  :  Instruction = "VOR.vv";
	    34'b1010111001010?100?????????????????  :  Instruction = "VOR.vx";
	    34'b1010111001010?011?????????????????  :  Instruction = "VOR.vi";
	    34'b1010111001011?000?????????????????  :  Instruction = "VXOR.vv";
	    34'b1010111001011?100?????????????????  :  Instruction = "VXOR.vx";
	    34'b1010111001011?011?????????????????  :  Instruction = "VXOR.vi";
	    34'b1010111010010?010?????????????????  :  Instruction = "VZEXT.vf2";
	    34'b1010111100101?000?????????????????  :  Instruction = "VSLL.vv";
	    34'b1010111100101?100?????????????????  :  Instruction = "VSLL.vx";
	    34'b1010111100101?011?????????????????  :  Instruction = "VSLL.vi";
	    34'b1010111101000?000?????????????????  :  Instruction = "VSRL.vv";
	    34'b1010111101000?100?????????????????  :  Instruction = "VSRL.vx";
	    34'b1010111101000?011?????????????????  :  Instruction = "VSRL.vi";
	    34'b1010111101001?000?????????????????  :  Instruction = "VSRA.vv";
	    34'b1010111101001?100?????????????????  :  Instruction = "VSRA.vx";
	    34'b1010111101001?011?????????????????  :  Instruction = "VSRA.vi";
	    34'b1010111101100?000?????????????????  :  Instruction = "VNSRL.wv";
	    34'b1010111101100?100?????????????????  :  Instruction = "VNSRL.wx";
	    34'b1010111101100?011?????????????????  :  Instruction = "VNSRL.wi";
	    34'b1010111101101?000?????????????????  :  Instruction = "VNSRA.wv";
	    34'b1010111101101?100?????????????????  :  Instruction = "VNSRA.wx";
	    34'b1010111101101?011?????????????????  :  Instruction = "VNSRA.wi";
	    34'b1010111011000?000?????????????????  :  Instruction = "VMSEQ.vv";
	    34'b1010111011000?100?????????????????  :  Instruction = "VMSEQ.vx";
	    34'b1010111011000?011?????????????????  :  Instruction = "VMSEQ.vi";
	    34'b1010111011001?000?????????????????  :  Instruction = "VMSNE.vv";
	    34'b1010111011001?100?????????????????  :  Instruction = "VMSNE.vx";
	    34'b1010111011001?011?????????????????  :  Instruction = "VMSNE.vi";
	    34'b1010111011010?000?????????????????  :  Instruction = "VMSLTU.vv";
	    34'b1010111011010?100?????????????????  :  Instruction = "VMSLTU.vx";
	    34'b1010111011011?000?????????????????  :  Instruction = "VMSLT.vv";
	    34'b1010111011011?100?????????????????  :  Instruction = "VMSLT.vx";
	    34'b1010111011100?000?????????????????  :  Instruction = "VMSLEU.vv";
	    34'b1010111011100?100?????????????????  :  Instruction = "VMSLEU.vx";
	    34'b1010111011100?011?????????????????  :  Instruction = "VMSLEU.vi";
	    34'b1010111011101?000?????????????????  :  Instruction = "VMSLE.vv";
	    34'b1010111011101?100?????????????????  :  Instruction = "VMSLE.vx";
	    34'b1010111011101?011?????????????????  :  Instruction = "VMSLE.vi";
	    34'b1010111011110?100?????????????????  :  Instruction = "VMSGTU.vx";
	    34'b1010111011110?011?????????????????  :  Instruction = "VMSGTU.vi";
	    34'b1010111011111?100?????????????????  :  Instruction = "VMSGT.vx";
	    34'b1010111011111?011?????????????????  :  Instruction = "VMSGT.vi";
	    34'b1010111000100?000?????????????????  :  Instruction = "VMINU.vv";
	    34'b1010111000100?100?????????????????  :  Instruction = "VMINU.vx";
	    34'b1010111000101?000?????????????????  :  Instruction = "VMIN.vv";
	    34'b1010111000101?100?????????????????  :  Instruction = "VMIN.vx";
	    34'b1010111000110?000?????????????????  :  Instruction = "VMAXU.vv";
	    34'b1010111000110?100?????????????????  :  Instruction = "VMAXU.vx";
	    34'b1010111000111?000?????????????????  :  Instruction = "VMAX.vv";
	    34'b1010111000111?100?????????????????  :  Instruction = "VMAX.vx";
	    34'b1010111100101?010?????????????????  :  Instruction = "VMUL.vv";
	    34'b1010111100101?110?????????????????  :  Instruction = "VMUL.vx";
	    34'b1010111100111?010?????????????????  :  Instruction = "VMULH.vv";
	    34'b1010111100111?110?????????????????  :  Instruction = "VMULH.vx";
	    34'b1010111100100?010?????????????????  :  Instruction = "VMULHU.vv";
	    34'b1010111100100?110?????????????????  :  Instruction = "VMULHU.vx";
	    34'b1010111100110?010?????????????????  :  Instruction = "VMULHSU.vv";
	    34'b1010111100110?110?????????????????  :  Instruction = "VMULHSU.vx";
	    34'b1010111111000?010?????????????????  :  Instruction = "VWMULU.vv";
	    34'b1010111111000?110?????????????????  :  Instruction = "VWMULU.vx";
	    34'b1010111111011?010?????????????????  :  Instruction = "VWMUL.vv";
	    34'b1010111111011?110?????????????????  :  Instruction = "VWMUL.vx";
	    34'b1010111111010?010?????????????????  :  Instruction = "VWMULSU.vv";
	    34'b1010111111010?110?????????????????  :  Instruction = "VWMULSU.vx";
	    34'b1010111101101?010?????????????????  :  Instruction = "VMACC.vv";
	    34'b1010111101101?110?????????????????  :  Instruction = "VMACC.vx";
	    34'b1010111101111?010?????????????????  :  Instruction = "VNMSAC.vv";
	    34'b1010111101111?110?????????????????  :  Instruction = "VNMSAC.vx";
	    34'b1010111101001?010?????????????????  :  Instruction = "VMADD.vv";
	    34'b1010111101001?110?????????????????  :  Instruction = "VMADD.vx";
	    34'b1010111101011?010?????????????????  :  Instruction = "VNMSUB.vv";
	    34'b1010111101011?110?????????????????  :  Instruction = "VNMSUB.vx";
	    34'b1010111111100?010?????????????????  :  Instruction = "VWMACCU.vv";
	    34'b1010111111100?110?????????????????  :  Instruction = "VWMACCU.vx";
	    34'b1010111111101?010?????????????????  :  Instruction = "VWMACC.vv";
	    34'b1010111111101?110?????????????????  :  Instruction = "VWMACC.vx";
	    34'b1010111111111?010?????????????????  :  Instruction = "VWMACCSU.vv";
	    34'b1010111111111?110?????????????????  :  Instruction = "VWMACCSU.vx";
	    34'b1010111111110?110?????????????????  :  Instruction = "VWMACCUS.vx";
	    34'b1010111010111?0000????????????????  :  Instruction = "VMERGE.vvm";
	    34'b1010111010111?1000????????????????  :  Instruction = "VMERGE.vxm";
	    34'b1010111010111?0110????????????????  :  Instruction = "VMERGE.vim";
	    34'b1010111010111?0001????????????????  :  Instruction = "VMV.v.v";
	    34'b1010111010111?1001????????????????  :  Instruction = "VMV.v.x";
	    34'b1010111010111?0111????????????????  :  Instruction = "VMV.v.i";
	    34'b1010111100000?000?????????????????  :  Instruction = "VSADDU.vv";
	    34'b1010111100000?100?????????????????  :  Instruction = "VSADDU.vx";
	    34'b1010111100000?011?????????????????  :  Instruction = "VSADDU.vi";
	    34'b1010111100001?000?????????????????  :  Instruction = "VSADD.vv";
	    34'b1010111100001?100?????????????????  :  Instruction = "VSADD.vx";
	    34'b1010111100001?011?????????????????  :  Instruction = "VSADD.vi";
	    34'b1010111100010?000?????????????????  :  Instruction = "VSSUBU.vv";
	    34'b1010111100010?100?????????????????  :  Instruction = "VSSUBU.vx";
	    34'b1010111100011?000?????????????????  :  Instruction = "VSSUB.vv";
	    34'b1010111100011?100?????????????????  :  Instruction = "VSSUB.vx";
	    34'b1010111001000?010?????????????????  :  Instruction = "VAADDU.vv";
	    34'b1010111001000?110?????????????????  :  Instruction = "VAADDU.vx";
	    34'b1010111001001?010?????????????????  :  Instruction = "VAADD.vv";
	    34'b1010111001001?110?????????????????  :  Instruction = "VAADD.vx";
	    34'b1010111001010?010?????????????????  :  Instruction = "VASUBU.vv";
	    34'b1010111001010?110?????????????????  :  Instruction = "VASUBU.vx";
	    34'b1010111001011?010?????????????????  :  Instruction = "VASUB.vv";
	    34'b1010111001011?110?????????????????  :  Instruction = "VASUB.vx";
	    34'b1010111100111?000?????????????????  :  Instruction = "VSMUL.vv";
	    34'b1010111100111?100?????????????????  :  Instruction = "VSMUL.vx";
	    34'b1010111100111?011?????????????????  :  Instruction = "VMV1R.v";
	    34'b1010111101010?000?????????????????  :  Instruction = "VSSRL.vv";
	    34'b1010111101010?100?????????????????  :  Instruction = "VSSRL.vx";
	    34'b1010111101010?011?????????????????  :  Instruction = "VSSRL.vi";
	    34'b1010111101011?000?????????????????  :  Instruction = "VSSRA.vv";
	    34'b1010111101011?100?????????????????  :  Instruction = "VSSRA.vx";
	    34'b1010111101011?011?????????????????  :  Instruction = "VSSRA.vi";
	    34'b1010111101110?000?????????????????  :  Instruction = "VNCLIPU.wv";
	    34'b1010111101110?100?????????????????  :  Instruction = "VNCLIPU.wx";
	    34'b1010111101110?011?????????????????  :  Instruction = "VNCLIPU.wi";
	    34'b1010111101111?000?????????????????  :  Instruction = "VNCLIP.wv";
	    34'b1010111101111?100?????????????????  :  Instruction = "VNCLIP.wx";
	    34'b1010111101111?011?????????????????  :  Instruction = "VNCLIP.wi";
	    34'b1010111000000?001?????????????????  :  Instruction = "VFADD.vv";
	    34'b1010111000000?101?????????????????  :  Instruction = "VFADD.vf";
	    34'b1010111000010?001?????????????????  :  Instruction = "VFSUB.vv";
	    34'b1010111000010?101?????????????????  :  Instruction = "VFSUB.vf";
	    34'b1010111100111?101?????????????????  :  Instruction = "VFRSUB.vf";
	    34'b1010111110000?001?????????????????  :  Instruction = "VFWADD.vv";
	    34'b1010111110000?101?????????????????  :  Instruction = "VFWADD.vf";
	    34'b1010111110100?001?????????????????  :  Instruction = "VFWADD.wv";
	    34'b1010111110100?101?????????????????  :  Instruction = "VFWADD.wf";
	    34'b1010111110010?001?????????????????  :  Instruction = "VFWSUB.vv";
	    34'b1010111110010?101?????????????????  :  Instruction = "VFWSUB.vf";
	    34'b1010111110110?001?????????????????  :  Instruction = "VFWSUB.wv";
	    34'b1010111110110?101?????????????????  :  Instruction = "VFWSUB.wf";
	    34'b1010111100100?001?????????????????  :  Instruction = "VFMUL.vv";
	    34'b1010111100100?101?????????????????  :  Instruction = "VFMUL.vf";
	    34'b1010111111000?001?????????????????  :  Instruction = "VFWMUL.vv";
	    34'b1010111111000?101?????????????????  :  Instruction = "VFWMUL.vf";
	    34'b1010111101100?001?????????????????  :  Instruction = "VFMACC.vv";
	    34'b1010111101100?101?????????????????  :  Instruction = "VFMACC.vf";
	    34'b1010111101101?001?????????????????  :  Instruction = "VFNMACC.vv";
	    34'b1010111101101?101?????????????????  :  Instruction = "VFNMACC.vf";
	    34'b1010111101110?001?????????????????  :  Instruction = "VFMSAC.vv";
	    34'b1010111101110?101?????????????????  :  Instruction = "VFMSAC.vf";
	    34'b1010111101111?001?????????????????  :  Instruction = "VFNMSAC.vv";
	    34'b1010111101111?101?????????????????  :  Instruction = "VFNMSAC.vf";
	    34'b1010111101000?001?????????????????  :  Instruction = "VFMADD.vv";
	    34'b1010111101000?101?????????????????  :  Instruction = "VFMADD.vf";
	    34'b1010111101001?001?????????????????  :  Instruction = "VFNMADD.vv";
	    34'b1010111101001?101?????????????????  :  Instruction = "VFNMADD.vf";
	    34'b1010111101010?001?????????????????  :  Instruction = "VFMSUB.vv";
	    34'b1010111101010?101?????????????????  :  Instruction = "VFMSUB.vf";
	    34'b1010111101011?001?????????????????  :  Instruction = "VFNMSUB.vv";
	    34'b1010111101011?101?????????????????  :  Instruction = "VFNMSUB.vf";
	    34'b1010111111100?001?????????????????  :  Instruction = "VFWMACC.vv";
	    34'b1010111111100?101?????????????????  :  Instruction = "VFWMACC.vf";
	    34'b1010111111101?001?????????????????  :  Instruction = "VFWNMACC.vv";
	    34'b1010111111101?101?????????????????  :  Instruction = "VFWNMACC.vf";
	    34'b1010111111110?001?????????????????  :  Instruction = "VFWMSAC.vv";
	    34'b1010111111110?101?????????????????  :  Instruction = "VFWMSAC.vf";
	    34'b1010111111111?001?????????????????  :  Instruction = "VFWNMSAC.vv";
	    34'b1010111111111?101?????????????????  :  Instruction = "VFWNMSAC.vf";
	    34'b1010111000100?001?????????????????  :  Instruction = "VFMIN.vv";
	    34'b1010111000100?101?????????????????  :  Instruction = "VFMIN.vf";
	    34'b1010111000110?001?????????????????  :  Instruction = "VFMAX.vv";
	    34'b1010111000110?101?????????????????  :  Instruction = "VFMAX.vf";
	    34'b1010111001000?001?????????????????  :  Instruction = "VFSGNJ.vv";
	    34'b1010111001000?101?????????????????  :  Instruction = "VFSGNJ.vf";
	    34'b1010111001001?001?????????????????  :  Instruction = "VFSGNJN.vv";
	    34'b1010111001001?101?????????????????  :  Instruction = "VFSGNJN.vf";
	    34'b1010111001010?001?????????????????  :  Instruction = "VFSGNJX.vv";
	    34'b1010111001010?101?????????????????  :  Instruction = "VFSGNJX.vf";
	    34'b1010111011000?001?????????????????  :  Instruction = "VMFEQ.vv";
	    34'b1010111011000?101?????????????????  :  Instruction = "VMFEQ.vf";
	    34'b1010111011100?001?????????????????  :  Instruction = "VMFNE.vv";
	    34'b1010111011100?101?????????????????  :  Instruction = "VMFNE.vf";
	    34'b1010111011011?001?????????????????  :  Instruction = "VMFLT.vv";
	    34'b1010111011011?101?????????????????  :  Instruction = "VMFLT.vf";
	    34'b1010111011001?001?????????????????  :  Instruction = "VMFLE.vv";
	    34'b1010111011001?101?????????????????  :  Instruction = "VMFLE.vf";
	    34'b1010111011101?101?????????????????  :  Instruction = "VMFGT.vf";
	    34'b1010111011111?101?????????????????  :  Instruction = "VMFGE.vf";
	    34'b1010111010011?001?????????????????  :  Instruction = "VFCLASS.v";
	    34'b1010111010111?101?????????????????  :  Instruction = "VFMERGE.vfm";
	    34'b1010111010111?1011????????????????  :  Instruction = "VFMV.v.f";
	    34'b1010111010010?001?????????????????  :  Instruction = "VFCVT.xu.f.v";
	    34'b1010111000000?010?????????????????  :  Instruction = "VREDSUM.vs";
	    34'b1010111000110?010?????????????????  :  Instruction = "VREDMAXU.vs";
	    34'b1010111000111?010?????????????????  :  Instruction = "VREDMAX.vs";
	    34'b1010111000100?010?????????????????  :  Instruction = "VREDMINU.vs";
	    34'b1010111000101?010?????????????????  :  Instruction = "VREDMIN.vs";
	    34'b1010111000001?010?????????????????  :  Instruction = "VREDAND.vs";
	    34'b1010111000010?010?????????????????  :  Instruction = "VREDOR.vs";
	    34'b1010111000011?010?????????????????  :  Instruction = "VREDXOR.vs";
	    34'b1010111110000?000?????????????????  :  Instruction = "VWREDSUMU.vs";
	    34'b1010111110001?000?????????????????  :  Instruction = "VWREDSUM.vs";
	    34'b1010111000011?001?????????????????  :  Instruction = "VFREDOSUM.vs";
	    34'b1010111000001?001?????????????????  :  Instruction = "VFREDSUM.vs";
	    34'b1010111000111?001?????????????????  :  Instruction = "VFREDMAX.vs";
	    34'b1010111000101?001?????????????????  :  Instruction = "VFREDMIN.vs";
	    34'b1010111110011?001?????????????????  :  Instruction = "VFWREDOSUM.vs";
	    34'b1010111110001?001?????????????????  :  Instruction = "VFWREDSUM.vs";
	    34'b1010111011001?010?????????????????  :  Instruction = "VMAND.mm";
	    34'b1010111011101?010?????????????????  :  Instruction = "VMNAND.mm";
	    34'b1010111011000?010?????????????????  :  Instruction = "VMANDNOT.mm";
	    34'b1010111011011?010?????????????????  :  Instruction = "VMXOR.mm";
	    34'b1010111011010?010?????????????????  :  Instruction = "VMOR.mm";
	    34'b1010111011110?010?????????????????  :  Instruction = "VMNOR.mm";
	    34'b1010111011100?010?????????????????  :  Instruction = "VMORNOT.mm";
	    34'b1010111011111?010?????????????????  :  Instruction = "VMXNOR.mm";
	    34'b1010111010000?010?????????????????  :  Instruction = "VPOPC.m";
	    34'b1010111010100?010?????????????????  :  Instruction = "VMSBF.m";
	    34'b1010111010000?110?????????????????  :  Instruction = "VMV.s.x";
	    34'b1010111010000?001?????????????????  :  Instruction = "VFMV.f.s";
	    34'b1010111010000?101?????????????????  :  Instruction = "VFMV.s.f";
	    34'b1010111001110?100?????????????????  :  Instruction = "VSLIDEUP.vx";
	    34'b1010111001110?011?????????????????  :  Instruction = "VSLIDEUP.vi";
	    34'b1010111001111?100?????????????????  :  Instruction = "VSLIDEDOWN.vx";
	    34'b1010111001111?011?????????????????  :  Instruction = "VSLIDEDOWN.vi";
	    34'b1010111001110?110?????????????????  :  Instruction = "VSLIDE1UP.vx";
	    34'b1010111001110?101?????????????????  :  Instruction = "VFSLIDE1UP.vf";
	    34'b1010111001111?110?????????????????  :  Instruction = "VSLIDE1DOWN.vx";
	    34'b1010111001111?101?????????????????  :  Instruction = "VFSLIDE1DOWN.vf";
	    34'b1010111001100?000?????????????????  :  Instruction = "VRGATHER.vv";
	    34'b1010111001100?100?????????????????  :  Instruction = "VRGATHER.vx";
	    34'b1010111001100?011?????????????????  :  Instruction = "VRGATHER.vi";
	    34'b1010111001110?000?????????????????  :  Instruction = "VRGATHEREI16.vv";
	    34'b1010111010111?010?????????????????  :  Instruction = "VCOMPRESS.vm";
	    34'b0000111???????000?00010100?0000???  :  Instruction = "vle8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000???  :  Instruction = "vle16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000???  :  Instruction = "vle32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000???  :  Instruction = "vle64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000???  :  Instruction = "vle8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000???  :  Instruction = "vle16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000???  :  Instruction = "vle32[ff].v,e8,mf4";
	    34'b0000111???????111?00011000?0000???  :  Instruction = "vle64[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000???  :  Instruction = "vle8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000???  :  Instruction = "vle16[ff].v,e8,mf2";
	    34'b0000111???????110?00011100?0000???  :  Instruction = "vle32[ff].v,e8,mf2";
	    34'b0000111???????111?00011100?0000???  :  Instruction = "vle64[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000???  :  Instruction = "vle8[ff].v,e8,m1";
	    34'b0000111???????101?00000000?0000???  :  Instruction = "vle16[ff].v,e8,m1";
	    34'b0000111???????110?00000000?0000???  :  Instruction = "vle32[ff].v,e8,m1";
	    34'b0000111???????111?00000000?0000???  :  Instruction = "vle64[ff].v,e8,m1";
	    34'b0000111???????000?00000100?0000???  :  Instruction = "vle8[ff].v,e8,m2";
	    34'b0000111???????101?00000100?0000???  :  Instruction = "vle16[ff].v,e8,m2";
	    34'b0000111???????110?00000100?0000???  :  Instruction = "vle32[ff].v,e8,m2";
	    34'b0000111???????000?00001000?0000???  :  Instruction = "vle8[ff].v,e8,m4";
	    34'b0000111???????101?00001000?0000???  :  Instruction = "vle16[ff].v,e8,m4";
	    34'b0000111???????000?00001100?0000???  :  Instruction = "vle8[ff].v,e8,m8";
	    34'b0000111???????000?000???0001000000  :  Instruction = "vl1re8.v,e8";
	    34'b0000111???????101?000???0001000000  :  Instruction = "vl1re16.v,e8";
	    34'b0000111???????110?000???0001000000  :  Instruction = "vl1re32.v,e8";
	    34'b0000111???????111?000???0001000000  :  Instruction = "vl1re64.v,e8";
	    34'b0000111???????000?00010110????????  :  Instruction = "vlse8.v,e8,mf8";
	    34'b0000111???????101?00010110????????  :  Instruction = "vlse16.v,e8,mf8";
	    34'b0000111???????110?00010110????????  :  Instruction = "vlse32.v,e8,mf8";
	    34'b0000111???????111?00010110????????  :  Instruction = "vlse64.v,e8,mf8";
	    34'b0000111???????000?00011010????????  :  Instruction = "vlse8.v,e8,mf4";
	    34'b0000111???????101?00011010????????  :  Instruction = "vlse16.v,e8,mf4";
	    34'b0000111???????110?00011010????????  :  Instruction = "vlse32.v,e8,mf4";
	    34'b0000111???????111?00011010????????  :  Instruction = "vlse64.v,e8,mf4";
	    34'b0000111???????000?00011110????????  :  Instruction = "vlse8.v,e8,mf2";
	    34'b0000111???????101?00011110????????  :  Instruction = "vlse16.v,e8,mf2";
	    34'b0000111???????110?00011110????????  :  Instruction = "vlse32.v,e8,mf2";
	    34'b0000111???????111?00011110????????  :  Instruction = "vlse64.v,e8,mf2";
	    34'b0000111???????000?00000010????????  :  Instruction = "vlse8.v,e8,m1";
	    34'b0000111???????101?00000010????????  :  Instruction = "vlse16.v,e8,m1";
	    34'b0000111???????110?00000010????????  :  Instruction = "vlse32.v,e8,m1";
	    34'b0000111???????111?00000010????????  :  Instruction = "vlse64.v,e8,m1";
	    34'b0000111???????000?00000110????????  :  Instruction = "vlse8.v,e8,m2";
	    34'b0000111???????101?00000110????????  :  Instruction = "vlse16.v,e8,m2";
	    34'b0000111???????110?00000110????????  :  Instruction = "vlse32.v,e8,m2";
	    34'b0000111???????000?00001010????????  :  Instruction = "vlse8.v,e8,m4";
	    34'b0000111???????101?00001010????????  :  Instruction = "vlse16.v,e8,m4";
	    34'b0000111???????000?00001110????????  :  Instruction = "vlse8.v,e8,m8";
	    34'b0000111???????000?000101?1????????  :  Instruction = "vl[uo]xei8.v,e8,mf8";
	    34'b0000111???????101?000101?1????????  :  Instruction = "vl[uo]xei16.v,e8,mf8";
	    34'b0000111???????110?000101?1????????  :  Instruction = "vl[uo]xei32.v,e8,mf8";
	    34'b0000111???????111?000101?1????????  :  Instruction = "vl[uo]xei64.v,e8,mf8";
	    34'b0000111???????000?000110?1????????  :  Instruction = "vl[uo]xei8.v,e8,mf4";
	    34'b0000111???????101?000110?1????????  :  Instruction = "vl[uo]xei16.v,e8,mf4";
	    34'b0000111???????110?000110?1????????  :  Instruction = "vl[uo]xei32.v,e8,mf4";
	    34'b0000111???????111?000110?1????????  :  Instruction = "vl[uo]xei64.v,e8,mf4";
	    34'b0000111???????000?000111?1????????  :  Instruction = "vl[uo]xei8.v,e8,mf2";
	    34'b0000111???????101?000111?1????????  :  Instruction = "vl[uo]xei16.v,e8,mf2";
	    34'b0000111???????110?000111?1????????  :  Instruction = "vl[uo]xei32.v,e8,mf2";
	    34'b0000111???????111?000111?1????????  :  Instruction = "vl[uo]xei64.v,e8,mf2";
	    34'b0000111???????000?000000?1????????  :  Instruction = "vl[uo]xei8.v,e8,m1";
	    34'b0000111???????101?000000?1????????  :  Instruction = "vl[uo]xei16.v,e8,m1";
	    34'b0000111???????110?000000?1????????  :  Instruction = "vl[uo]xei32.v,e8,m1";
	    34'b0000111???????111?000000?1????????  :  Instruction = "vl[uo]xei64.v,e8,m1";
	    34'b0000111???????000?000001?1????????  :  Instruction = "vl[uo]xei8.v,e8,m2";
	    34'b0000111???????101?000001?1????????  :  Instruction = "vl[uo]xei16.v,e8,m2";
	    34'b0000111???????110?000001?1????????  :  Instruction = "vl[uo]xei32.v,e8,m2";
	    34'b0000111???????000?000010?1????????  :  Instruction = "vl[uo]xei8.v,e8,m4";
	    34'b0000111???????101?000010?1????????  :  Instruction = "vl[uo]xei16.v,e8,m4";
	    34'b0000111???????000?000011?1????????  :  Instruction = "vl[uo]xei8.v,e8,m8";
	    34'b0000111???????000?00010100?0000001  :  Instruction = "vlseg2e8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000001  :  Instruction = "vlseg2e16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000001  :  Instruction = "vlseg2e32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000001  :  Instruction = "vlseg2e64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000001  :  Instruction = "vlseg2e8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000001  :  Instruction = "vlseg2e16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000001  :  Instruction = "vlseg2e32[ff].v,e8,mf4";
	    34'b0000111???????111?00011000?0000001  :  Instruction = "vlseg2e64[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000001  :  Instruction = "vlseg2e8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000001  :  Instruction = "vlseg2e16[ff].v,e8,mf2";
	    34'b0000111???????110?00011100?0000001  :  Instruction = "vlseg2e32[ff].v,e8,mf2";
	    34'b0000111???????111?00011100?0000001  :  Instruction = "vlseg2e64[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000001  :  Instruction = "vlseg2e8[ff].v,e8,m1";
	    34'b0000111???????101?00000000?0000001  :  Instruction = "vlseg2e16[ff].v,e8,m1";
	    34'b0000111???????110?00000000?0000001  :  Instruction = "vlseg2e32[ff].v,e8,m1";
	    34'b0000111???????000?00000100?0000001  :  Instruction = "vlseg2e8[ff].v,e8,m2";
	    34'b0000111???????101?00000100?0000001  :  Instruction = "vlseg2e16[ff].v,e8,m2";
	    34'b0000111???????000?00001000?0000001  :  Instruction = "vlseg2e8[ff].v,e8,m4";
	    34'b0000111???????111?00001100?0000001  :  Instruction = "vlseg2e64[ff].v,e8,m8";
	    34'b0000111???????000?000???0001000001  :  Instruction = "vl2re8.v,e8";
	    34'b0000111???????101?000???0001000001  :  Instruction = "vl2re16.v,e8";
	    34'b0000111???????110?000???0001000001  :  Instruction = "vl2re32.v,e8";
	    34'b0000111???????111?000???0001000001  :  Instruction = "vl2re64.v,e8";
	    34'b0000111???????000?00010110?????001  :  Instruction = "vlsseg2e8.v,e8,mf8";
	    34'b0000111???????101?00010110?????001  :  Instruction = "vlsseg2e16.v,e8,mf8";
	    34'b0000111???????110?00010110?????001  :  Instruction = "vlsseg2e32.v,e8,mf8";
	    34'b0000111???????111?00010110?????001  :  Instruction = "vlsseg2e64.v,e8,mf8";
	    34'b0000111???????000?00011010?????001  :  Instruction = "vlsseg2e8.v,e8,mf4";
	    34'b0000111???????101?00011010?????001  :  Instruction = "vlsseg2e16.v,e8,mf4";
	    34'b0000111???????110?00011010?????001  :  Instruction = "vlsseg2e32.v,e8,mf4";
	    34'b0000111???????111?00011010?????001  :  Instruction = "vlsseg2e64.v,e8,mf4";
	    34'b0000111???????000?00011110?????001  :  Instruction = "vlsseg2e8.v,e8,mf2";
	    34'b0000111???????101?00011110?????001  :  Instruction = "vlsseg2e16.v,e8,mf2";
	    34'b0000111???????110?00011110?????001  :  Instruction = "vlsseg2e32.v,e8,mf2";
	    34'b0000111???????111?00011110?????001  :  Instruction = "vlsseg2e64.v,e8,mf2";
	    34'b0000111???????000?00000010?????001  :  Instruction = "vlsseg2e8.v,e8,m1";
	    34'b0000111???????101?00000010?????001  :  Instruction = "vlsseg2e16.v,e8,m1";
	    34'b0000111???????110?00000010?????001  :  Instruction = "vlsseg2e32.v,e8,m1";
	    34'b0000111???????000?00000110?????001  :  Instruction = "vlsseg2e8.v,e8,m2";
	    34'b0000111???????101?00000110?????001  :  Instruction = "vlsseg2e16.v,e8,m2";
	    34'b0000111???????000?00001010?????001  :  Instruction = "vlsseg2e8.v,e8,m4";
	    34'b0000111???????000?000101?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e8,mf8";
	    34'b0000111???????101?000101?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e8,mf8";
	    34'b0000111???????110?000101?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e8,mf8";
	    34'b0000111???????111?000101?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e8,mf8";
	    34'b0000111???????000?000110?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e8,mf4";
	    34'b0000111???????101?000110?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e8,mf4";
	    34'b0000111???????110?000110?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e8,mf4";
	    34'b0000111???????111?000110?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e8,mf4";
	    34'b0000111???????000?000111?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e8,mf2";
	    34'b0000111???????101?000111?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e8,mf2";
	    34'b0000111???????110?000111?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e8,mf2";
	    34'b0000111???????111?000111?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e8,mf2";
	    34'b0000111???????000?000000?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e8,m1";
	    34'b0000111???????101?000000?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e8,m1";
	    34'b0000111???????110?000000?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e8,m1";
	    34'b0000111???????111?000000?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e8,m1";
	    34'b0000111???????000?000001?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e8,m2";
	    34'b0000111???????101?000001?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e8,m2";
	    34'b0000111???????110?000001?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e8,m2";
	    34'b0000111???????000?000010?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e8,m4";
	    34'b0000111???????101?000010?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e8,m4";
	    34'b0000111???????000?00010100?0000010  :  Instruction = "vlseg3e8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000010  :  Instruction = "vlseg3e16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000010  :  Instruction = "vlseg3e32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000010  :  Instruction = "vlseg3e64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000010  :  Instruction = "vlseg3e8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000010  :  Instruction = "vlseg3e16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000010  :  Instruction = "vlseg3e32[ff].v,e8,mf4";
	    34'b0000111???????111?00011000?0000010  :  Instruction = "vlseg3e64[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000010  :  Instruction = "vlseg3e8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000010  :  Instruction = "vlseg3e16[ff].v,e8,mf2";
	    34'b0000111???????110?00011100?0000010  :  Instruction = "vlseg3e32[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000010  :  Instruction = "vlseg3e8[ff].v,e8,m1";
	    34'b0000111???????101?00000000?0000010  :  Instruction = "vlseg3e16[ff].v,e8,m1";
	    34'b0000111???????000?00000100?0000010  :  Instruction = "vlseg3e8[ff].v,e8,m2";
	    34'b0000111???????000?00010110?????010  :  Instruction = "vlsseg3e8.v,e8,mf8";
	    34'b0000111???????101?00010110?????010  :  Instruction = "vlsseg3e16.v,e8,mf8";
	    34'b0000111???????110?00010110?????010  :  Instruction = "vlsseg3e32.v,e8,mf8";
	    34'b0000111???????111?00010110?????010  :  Instruction = "vlsseg3e64.v,e8,mf8";
	    34'b0000111???????000?00011010?????010  :  Instruction = "vlsseg3e8.v,e8,mf4";
	    34'b0000111???????101?00011010?????010  :  Instruction = "vlsseg3e16.v,e8,mf4";
	    34'b0000111???????110?00011010?????010  :  Instruction = "vlsseg3e32.v,e8,mf4";
	    34'b0000111???????111?00011010?????010  :  Instruction = "vlsseg3e64.v,e8,mf4";
	    34'b0000111???????000?00011110?????010  :  Instruction = "vlsseg3e8.v,e8,mf2";
	    34'b0000111???????101?00011110?????010  :  Instruction = "vlsseg3e16.v,e8,mf2";
	    34'b0000111???????110?00011110?????010  :  Instruction = "vlsseg3e32.v,e8,mf2";
	    34'b0000111???????000?00000010?????010  :  Instruction = "vlsseg3e8.v,e8,m1";
	    34'b0000111???????101?00000010?????010  :  Instruction = "vlsseg3e16.v,e8,m1";
	    34'b0000111???????000?00000110?????010  :  Instruction = "vlsseg3e8.v,e8,m2";
	    34'b0000111???????000?000101?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e8,mf8";
	    34'b0000111???????101?000101?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e8,mf8";
	    34'b0000111???????110?000101?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e8,mf8";
	    34'b0000111???????111?000101?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e8,mf8";
	    34'b0000111???????000?000110?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e8,mf4";
	    34'b0000111???????101?000110?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e8,mf4";
	    34'b0000111???????110?000110?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e8,mf4";
	    34'b0000111???????111?000110?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e8,mf4";
	    34'b0000111???????000?000111?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e8,mf2";
	    34'b0000111???????101?000111?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e8,mf2";
	    34'b0000111???????110?000111?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e8,mf2";
	    34'b0000111???????111?000111?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e8,mf2";
	    34'b0000111???????000?000000?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e8,m1";
	    34'b0000111???????101?000000?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e8,m1";
	    34'b0000111???????110?000000?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e8,m1";
	    34'b0000111???????111?000000?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e8,m1";
	    34'b0000111???????000?000001?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e8,m2";
	    34'b0000111???????101?000001?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e8,m2";
	    34'b0000111???????110?000001?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e8,m2";
	    34'b0000111???????000?00010100?0000011  :  Instruction = "vlseg4e8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000011  :  Instruction = "vlseg4e16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000011  :  Instruction = "vlseg4e32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000011  :  Instruction = "vlseg4e64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000011  :  Instruction = "vlseg4e8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000011  :  Instruction = "vlseg4e16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000011  :  Instruction = "vlseg4e32[ff].v,e8,mf4";
	    34'b0000111???????111?00011000?0000011  :  Instruction = "vlseg4e64[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000011  :  Instruction = "vlseg4e8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000011  :  Instruction = "vlseg4e16[ff].v,e8,mf2";
	    34'b0000111???????110?00011100?0000011  :  Instruction = "vlseg4e32[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000011  :  Instruction = "vlseg4e8[ff].v,e8,m1";
	    34'b0000111???????101?00000000?0000011  :  Instruction = "vlseg4e16[ff].v,e8,m1";
	    34'b0000111???????000?00000100?0000011  :  Instruction = "vlseg4e8[ff].v,e8,m2";
	    34'b0000111???????000?00010110?????011  :  Instruction = "vlsseg4e8.v,e8,mf8";
	    34'b0000111???????101?00010110?????011  :  Instruction = "vlsseg4e16.v,e8,mf8";
	    34'b0000111???????110?00010110?????011  :  Instruction = "vlsseg4e32.v,e8,mf8";
	    34'b0000111???????111?00010110?????011  :  Instruction = "vlsseg4e64.v,e8,mf8";
	    34'b0000111???????000?00011010?????011  :  Instruction = "vlsseg4e8.v,e8,mf4";
	    34'b0000111???????101?00011010?????011  :  Instruction = "vlsseg4e16.v,e8,mf4";
	    34'b0000111???????110?00011010?????011  :  Instruction = "vlsseg4e32.v,e8,mf4";
	    34'b0000111???????111?00011010?????011  :  Instruction = "vlsseg4e64.v,e8,mf4";
	    34'b0000111???????000?00011110?????011  :  Instruction = "vlsseg4e8.v,e8,mf2";
	    34'b0000111???????101?00011110?????011  :  Instruction = "vlsseg4e16.v,e8,mf2";
	    34'b0000111???????110?00011110?????011  :  Instruction = "vlsseg4e32.v,e8,mf2";
	    34'b0000111???????000?00000010?????011  :  Instruction = "vlsseg4e8.v,e8,m1";
	    34'b0000111???????101?00000010?????011  :  Instruction = "vlsseg4e16.v,e8,m1";
	    34'b0000111???????000?00000110?????011  :  Instruction = "vlsseg4e8.v,e8,m2";
	    34'b0000111???????000?000???0001000011  :  Instruction = "vl4re8.v,e8";
	    34'b0000111???????101?000???0001000011  :  Instruction = "vl4re16.v,e8";
	    34'b0000111???????110?000???0001000011  :  Instruction = "vl4re32.v,e8";
	    34'b0000111???????111?000???0001000011  :  Instruction = "vl4re64.v,e8";
	    34'b0000111???????000?000101?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e8,mf8";
	    34'b0000111???????101?000101?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e8,mf8";
	    34'b0000111???????110?000101?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e8,mf8";
	    34'b0000111???????111?000101?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e8,mf8";
	    34'b0000111???????000?000110?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e8,mf4";
	    34'b0000111???????101?000110?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e8,mf4";
	    34'b0000111???????110?000110?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e8,mf4";
	    34'b0000111???????111?000110?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e8,mf4";
	    34'b0000111???????000?000111?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e8,mf2";
	    34'b0000111???????101?000111?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e8,mf2";
	    34'b0000111???????110?000111?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e8,mf2";
	    34'b0000111???????111?000111?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e8,mf2";
	    34'b0000111???????000?000000?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e8,m1";
	    34'b0000111???????101?000000?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e8,m1";
	    34'b0000111???????110?000000?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e8,m1";
	    34'b0000111???????111?000000?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e8,m1";
	    34'b0000111???????000?000001?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e8,m2";
	    34'b0000111???????101?000001?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e8,m2";
	    34'b0000111???????110?000001?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e8,m2";
	    34'b0000111???????000?00010100?0000100  :  Instruction = "vlseg5e8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000100  :  Instruction = "vlseg5e16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000100  :  Instruction = "vlseg5e32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000100  :  Instruction = "vlseg5e64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000100  :  Instruction = "vlseg5e8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000100  :  Instruction = "vlseg5e16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000100  :  Instruction = "vlseg5e32[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000100  :  Instruction = "vlseg5e8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000100  :  Instruction = "vlseg5e16[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000100  :  Instruction = "vlseg5e8[ff].v,e8,m1";
	    34'b0000111???????000?00010110?????100  :  Instruction = "vlsseg5e8.v,e8,mf8";
	    34'b0000111???????101?00010110?????100  :  Instruction = "vlsseg5e16.v,e8,mf8";
	    34'b0000111???????110?00010110?????100  :  Instruction = "vlsseg5e32.v,e8,mf8";
	    34'b0000111???????111?00010110?????100  :  Instruction = "vlsseg5e64.v,e8,mf8";
	    34'b0000111???????000?00011010?????100  :  Instruction = "vlsseg5e8.v,e8,mf4";
	    34'b0000111???????101?00011010?????100  :  Instruction = "vlsseg5e16.v,e8,mf4";
	    34'b0000111???????110?00011010?????100  :  Instruction = "vlsseg5e32.v,e8,mf4";
	    34'b0000111???????000?00011110?????100  :  Instruction = "vlsseg5e8.v,e8,mf2";
	    34'b0000111???????101?00011110?????100  :  Instruction = "vlsseg5e16.v,e8,mf2";
	    34'b0000111???????000?00000010?????100  :  Instruction = "vlsseg5e8.v,e8,m1";
	    34'b0000111???????000?000101?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e8,mf8";
	    34'b0000111???????101?000101?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e8,mf8";
	    34'b0000111???????110?000101?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e8,mf8";
	    34'b0000111???????111?000101?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e8,mf8";
	    34'b0000111???????000?000110?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e8,mf4";
	    34'b0000111???????101?000110?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e8,mf4";
	    34'b0000111???????110?000110?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e8,mf4";
	    34'b0000111???????111?000110?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e8,mf4";
	    34'b0000111???????000?000111?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e8,mf2";
	    34'b0000111???????101?000111?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e8,mf2";
	    34'b0000111???????110?000111?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e8,mf2";
	    34'b0000111???????111?000111?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e8,mf2";
	    34'b0000111???????000?000000?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e8,m1";
	    34'b0000111???????101?000000?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e8,m1";
	    34'b0000111???????110?000000?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e8,m1";
	    34'b0000111???????111?000000?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e8,m1";
	    34'b0000111???????000?00010100?0000101  :  Instruction = "vlseg6e8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000101  :  Instruction = "vlseg6e16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000101  :  Instruction = "vlseg6e32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000101  :  Instruction = "vlseg6e64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000101  :  Instruction = "vlseg6e8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000101  :  Instruction = "vlseg6e16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000101  :  Instruction = "vlseg6e32[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000101  :  Instruction = "vlseg6e8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000101  :  Instruction = "vlseg6e16[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000101  :  Instruction = "vlseg6e8[ff].v,e8,m1";
	    34'b0000111???????000?00010110?????101  :  Instruction = "vlsseg6e8.v,e8,mf8";
	    34'b0000111???????101?00010110?????101  :  Instruction = "vlsseg6e16.v,e8,mf8";
	    34'b0000111???????110?00010110?????101  :  Instruction = "vlsseg6e32.v,e8,mf8";
	    34'b0000111???????111?00010110?????101  :  Instruction = "vlsseg6e64.v,e8,mf8";
	    34'b0000111???????000?00011010?????101  :  Instruction = "vlsseg6e8.v,e8,mf4";
	    34'b0000111???????101?00011010?????101  :  Instruction = "vlsseg6e16.v,e8,mf4";
	    34'b0000111???????110?00011010?????101  :  Instruction = "vlsseg6e32.v,e8,mf4";
	    34'b0000111???????000?00011110?????101  :  Instruction = "vlsseg6e8.v,e8,mf2";
	    34'b0000111???????101?00011110?????101  :  Instruction = "vlsseg6e16.v,e8,mf2";
	    34'b0000111???????000?00000010?????101  :  Instruction = "vlsseg6e8.v,e8,m1";
	    34'b0000111???????000?000101?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e8,mf8";
	    34'b0000111???????101?000101?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e8,mf8";
	    34'b0000111???????110?000101?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e8,mf8";
	    34'b0000111???????111?000101?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e8,mf8";
	    34'b0000111???????000?000110?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e8,mf4";
	    34'b0000111???????101?000110?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e8,mf4";
	    34'b0000111???????110?000110?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e8,mf4";
	    34'b0000111???????111?000110?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e8,mf4";
	    34'b0000111???????000?000111?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e8,mf2";
	    34'b0000111???????101?000111?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e8,mf2";
	    34'b0000111???????110?000111?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e8,mf2";
	    34'b0000111???????111?000111?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e8,mf2";
	    34'b0000111???????000?000000?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e8,m1";
	    34'b0000111???????101?000000?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e8,m1";
	    34'b0000111???????110?000000?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e8,m1";
	    34'b0000111???????111?000000?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e8,m1";
	    34'b0000111???????000?00010100?0000110  :  Instruction = "vlseg7e8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000110  :  Instruction = "vlseg7e16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000110  :  Instruction = "vlseg7e32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000110  :  Instruction = "vlseg7e64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000110  :  Instruction = "vlseg7e8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000110  :  Instruction = "vlseg7e16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000110  :  Instruction = "vlseg7e32[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000110  :  Instruction = "vlseg7e8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000110  :  Instruction = "vlseg7e16[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000110  :  Instruction = "vlseg7e8[ff].v,e8,m1";
	    34'b0000111???????000?00010110?????110  :  Instruction = "vlsseg7e8.v,e8,mf8";
	    34'b0000111???????101?00010110?????110  :  Instruction = "vlsseg7e16.v,e8,mf8";
	    34'b0000111???????110?00010110?????110  :  Instruction = "vlsseg7e32.v,e8,mf8";
	    34'b0000111???????111?00010110?????110  :  Instruction = "vlsseg7e64.v,e8,mf8";
	    34'b0000111???????000?00011010?????110  :  Instruction = "vlsseg7e8.v,e8,mf4";
	    34'b0000111???????101?00011010?????110  :  Instruction = "vlsseg7e16.v,e8,mf4";
	    34'b0000111???????110?00011010?????110  :  Instruction = "vlsseg7e32.v,e8,mf4";
	    34'b0000111???????000?00011110?????110  :  Instruction = "vlsseg7e8.v,e8,mf2";
	    34'b0000111???????101?00011110?????110  :  Instruction = "vlsseg7e16.v,e8,mf2";
	    34'b0000111???????000?00000010?????110  :  Instruction = "vlsseg7e8.v,e8,m1";
	    34'b0000111???????000?000101?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e8,mf8";
	    34'b0000111???????101?000101?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e8,mf8";
	    34'b0000111???????110?000101?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e8,mf8";
	    34'b0000111???????111?000101?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e8,mf8";
	    34'b0000111???????000?000110?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e8,mf4";
	    34'b0000111???????101?000110?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e8,mf4";
	    34'b0000111???????110?000110?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e8,mf4";
	    34'b0000111???????111?000110?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e8,mf4";
	    34'b0000111???????000?000111?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e8,mf2";
	    34'b0000111???????101?000111?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e8,mf2";
	    34'b0000111???????110?000111?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e8,mf2";
	    34'b0000111???????111?000111?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e8,mf2";
	    34'b0000111???????000?000000?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e8,m1";
	    34'b0000111???????101?000000?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e8,m1";
	    34'b0000111???????110?000000?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e8,m1";
	    34'b0000111???????111?000000?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e8,m1";
	    34'b0000111???????000?00010100?0000111  :  Instruction = "vlseg8e8[ff].v,e8,mf8";
	    34'b0000111???????101?00010100?0000111  :  Instruction = "vlseg8e16[ff].v,e8,mf8";
	    34'b0000111???????110?00010100?0000111  :  Instruction = "vlseg8e32[ff].v,e8,mf8";
	    34'b0000111???????111?00010100?0000111  :  Instruction = "vlseg8e64[ff].v,e8,mf8";
	    34'b0000111???????000?00011000?0000111  :  Instruction = "vlseg8e8[ff].v,e8,mf4";
	    34'b0000111???????101?00011000?0000111  :  Instruction = "vlseg8e16[ff].v,e8,mf4";
	    34'b0000111???????110?00011000?0000111  :  Instruction = "vlseg8e32[ff].v,e8,mf4";
	    34'b0000111???????000?00011100?0000111  :  Instruction = "vlseg8e8[ff].v,e8,mf2";
	    34'b0000111???????101?00011100?0000111  :  Instruction = "vlseg8e16[ff].v,e8,mf2";
	    34'b0000111???????000?00000000?0000111  :  Instruction = "vlseg8e8[ff].v,e8,m1";
	    34'b0000111???????000?000???0001000111  :  Instruction = "vl8re8.v,e8";
	    34'b0000111???????101?000???0001000111  :  Instruction = "vl8re16.v,e8";
	    34'b0000111???????110?000???0001000111  :  Instruction = "vl8re32.v,e8";
	    34'b0000111???????111?000???0001000111  :  Instruction = "vl8re64.v,e8";
	    34'b0000111???????000?00010110?????111  :  Instruction = "vlsseg8e8.v,e8,mf8";
	    34'b0000111???????101?00010110?????111  :  Instruction = "vlsseg8e16.v,e8,mf8";
	    34'b0000111???????110?00010110?????111  :  Instruction = "vlsseg8e32.v,e8,mf8";
	    34'b0000111???????111?00010110?????111  :  Instruction = "vlsseg8e64.v,e8,mf8";
	    34'b0000111???????000?00011010?????111  :  Instruction = "vlsseg8e8.v,e8,mf4";
	    34'b0000111???????101?00011010?????111  :  Instruction = "vlsseg8e16.v,e8,mf4";
	    34'b0000111???????110?00011010?????111  :  Instruction = "vlsseg8e32.v,e8,mf4";
	    34'b0000111???????000?00011110?????111  :  Instruction = "vlsseg8e8.v,e8,mf2";
	    34'b0000111???????101?00011110?????111  :  Instruction = "vlsseg8e16.v,e8,mf2";
	    34'b0000111???????000?00000010?????111  :  Instruction = "vlsseg8e8.v,e8,m1";
	    34'b0000111???????000?000101?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e8,mf8";
	    34'b0000111???????101?000101?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e8,mf8";
	    34'b0000111???????110?000101?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e8,mf8";
	    34'b0000111???????111?000101?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e8,mf8";
	    34'b0000111???????000?000110?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e8,mf4";
	    34'b0000111???????101?000110?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e8,mf4";
	    34'b0000111???????110?000110?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e8,mf4";
	    34'b0000111???????111?000110?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e8,mf4";
	    34'b0000111???????000?000111?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e8,mf2";
	    34'b0000111???????101?000111?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e8,mf2";
	    34'b0000111???????110?000111?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e8,mf2";
	    34'b0000111???????111?000111?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e8,mf2";
	    34'b0000111???????000?000000?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e8,m1";
	    34'b0000111???????101?000000?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e8,m1";
	    34'b0000111???????110?000000?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e8,m1";
	    34'b0000111???????111?000000?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e8,m1";
	    34'b0100111???????000?00010100?0000???  :  Instruction = "vse8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000???  :  Instruction = "vse16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000???  :  Instruction = "vse32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000???  :  Instruction = "vse64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000???  :  Instruction = "vse8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000???  :  Instruction = "vse16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000???  :  Instruction = "vse32[ff].v,e8,mf4";
	    34'b0100111???????111?00011000?0000???  :  Instruction = "vse64[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000???  :  Instruction = "vse8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000???  :  Instruction = "vse16[ff].v,e8,mf2";
	    34'b0100111???????110?00011100?0000???  :  Instruction = "vse32[ff].v,e8,mf2";
	    34'b0100111???????111?00011100?0000???  :  Instruction = "vse64[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000???  :  Instruction = "vse8[ff].v,e8,m1";
	    34'b0100111???????101?00000000?0000???  :  Instruction = "vse16[ff].v,e8,m1";
	    34'b0100111???????110?00000000?0000???  :  Instruction = "vse32[ff].v,e8,m1";
	    34'b0100111???????111?00000000?0000???  :  Instruction = "vse64[ff].v,e8,m1";
	    34'b0100111???????000?00000100?0000???  :  Instruction = "vse8[ff].v,e8,m2";
	    34'b0100111???????101?00000100?0000???  :  Instruction = "vse16[ff].v,e8,m2";
	    34'b0100111???????110?00000100?0000???  :  Instruction = "vse32[ff].v,e8,m2";
	    34'b0100111???????000?00001000?0000???  :  Instruction = "vse8[ff].v,e8,m4";
	    34'b0100111???????101?00001000?0000???  :  Instruction = "vse16[ff].v,e8,m4";
	    34'b0100111???????000?00001100?0000???  :  Instruction = "vse8[ff].v,e8,m8";
	    34'b0100111???????000?000???0001000000  :  Instruction = "vs1r.v,e8";
	    34'b0100111???????000?00010110????????  :  Instruction = "vsse8.v,e8,mf8";
	    34'b0100111???????101?00010110????????  :  Instruction = "vsse16.v,e8,mf8";
	    34'b0100111???????110?00010110????????  :  Instruction = "vsse32.v,e8,mf8";
	    34'b0100111???????111?00010110????????  :  Instruction = "vsse64.v,e8,mf8";
	    34'b0100111???????000?00011010????????  :  Instruction = "vsse8.v,e8,mf4";
	    34'b0100111???????101?00011010????????  :  Instruction = "vsse16.v,e8,mf4";
	    34'b0100111???????110?00011010????????  :  Instruction = "vsse32.v,e8,mf4";
	    34'b0100111???????111?00011010????????  :  Instruction = "vsse64.v,e8,mf4";
	    34'b0100111???????000?00011110????????  :  Instruction = "vsse8.v,e8,mf2";
	    34'b0100111???????101?00011110????????  :  Instruction = "vsse16.v,e8,mf2";
	    34'b0100111???????110?00011110????????  :  Instruction = "vsse32.v,e8,mf2";
	    34'b0100111???????111?00011110????????  :  Instruction = "vsse64.v,e8,mf2";
	    34'b0100111???????000?00000010????????  :  Instruction = "vsse8.v,e8,m1";
	    34'b0100111???????101?00000010????????  :  Instruction = "vsse16.v,e8,m1";
	    34'b0100111???????110?00000010????????  :  Instruction = "vsse32.v,e8,m1";
	    34'b0100111???????111?00000010????????  :  Instruction = "vsse64.v,e8,m1";
	    34'b0100111???????000?00000110????????  :  Instruction = "vsse8.v,e8,m2";
	    34'b0100111???????101?00000110????????  :  Instruction = "vsse16.v,e8,m2";
	    34'b0100111???????110?00000110????????  :  Instruction = "vsse32.v,e8,m2";
	    34'b0100111???????000?00001010????????  :  Instruction = "vsse8.v,e8,m4";
	    34'b0100111???????101?00001010????????  :  Instruction = "vsse16.v,e8,m4";
	    34'b0100111???????000?00001110????????  :  Instruction = "vsse8.v,e8,m8";
	    34'b0100111???????000?000101?1????????  :  Instruction = "vs[uo]xei8.v,e8,mf8";
	    34'b0100111???????101?000101?1????????  :  Instruction = "vs[uo]xei16.v,e8,mf8";
	    34'b0100111???????110?000101?1????????  :  Instruction = "vs[uo]xei32.v,e8,mf8";
	    34'b0100111???????111?000101?1????????  :  Instruction = "vs[uo]xei64.v,e8,mf8";
	    34'b0100111???????000?000110?1????????  :  Instruction = "vs[uo]xei8.v,e8,mf4";
	    34'b0100111???????101?000110?1????????  :  Instruction = "vs[uo]xei16.v,e8,mf4";
	    34'b0100111???????110?000110?1????????  :  Instruction = "vs[uo]xei32.v,e8,mf4";
	    34'b0100111???????111?000110?1????????  :  Instruction = "vs[uo]xei64.v,e8,mf4";
	    34'b0100111???????000?000111?1????????  :  Instruction = "vs[uo]xei8.v,e8,mf2";
	    34'b0100111???????101?000111?1????????  :  Instruction = "vs[uo]xei16.v,e8,mf2";
	    34'b0100111???????110?000111?1????????  :  Instruction = "vs[uo]xei32.v,e8,mf2";
	    34'b0100111???????111?000111?1????????  :  Instruction = "vs[uo]xei64.v,e8,mf2";
	    34'b0100111???????000?000000?1????????  :  Instruction = "vs[uo]xei8.v,e8,m1";
	    34'b0100111???????101?000000?1????????  :  Instruction = "vs[uo]xei16.v,e8,m1";
	    34'b0100111???????110?000000?1????????  :  Instruction = "vs[uo]xei32.v,e8,m1";
	    34'b0100111???????111?000000?1????????  :  Instruction = "vs[uo]xei64.v,e8,m1";
	    34'b0100111???????000?000001?1????????  :  Instruction = "vs[uo]xei8.v,e8,m2";
	    34'b0100111???????101?000001?1????????  :  Instruction = "vs[uo]xei16.v,e8,m2";
	    34'b0100111???????110?000001?1????????  :  Instruction = "vs[uo]xei32.v,e8,m2";
	    34'b0100111???????000?000010?1????????  :  Instruction = "vs[uo]xei8.v,e8,m4";
	    34'b0100111???????101?000010?1????????  :  Instruction = "vs[uo]xei16.v,e8,m4";
	    34'b0100111???????000?000011?1????????  :  Instruction = "vs[uo]xei8.v,e8,m8";
	    34'b0100111???????000?00010100?0000001  :  Instruction = "vsseg2e8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000001  :  Instruction = "vsseg2e16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000001  :  Instruction = "vsseg2e32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000001  :  Instruction = "vsseg2e64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000001  :  Instruction = "vsseg2e8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000001  :  Instruction = "vsseg2e16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000001  :  Instruction = "vsseg2e32[ff].v,e8,mf4";
	    34'b0100111???????111?00011000?0000001  :  Instruction = "vsseg2e64[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000001  :  Instruction = "vsseg2e8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000001  :  Instruction = "vsseg2e16[ff].v,e8,mf2";
	    34'b0100111???????110?00011100?0000001  :  Instruction = "vsseg2e32[ff].v,e8,mf2";
	    34'b0100111???????111?00011100?0000001  :  Instruction = "vsseg2e64[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000001  :  Instruction = "vsseg2e8[ff].v,e8,m1";
	    34'b0100111???????101?00000000?0000001  :  Instruction = "vsseg2e16[ff].v,e8,m1";
	    34'b0100111???????110?00000000?0000001  :  Instruction = "vsseg2e32[ff].v,e8,m1";
	    34'b0100111???????000?00000100?0000001  :  Instruction = "vsseg2e8[ff].v,e8,m2";
	    34'b0100111???????101?00000100?0000001  :  Instruction = "vsseg2e16[ff].v,e8,m2";
	    34'b0100111???????000?00001000?0000001  :  Instruction = "vsseg2e8[ff].v,e8,m4";
	    34'b0100111???????000?000???0001000001  :  Instruction = "vs2r.v,e8";
	    34'b0100111???????000?00010110?????001  :  Instruction = "vssseg2e8.v,e8,mf8";
	    34'b0100111???????101?00010110?????001  :  Instruction = "vssseg2e16.v,e8,mf8";
	    34'b0100111???????110?00010110?????001  :  Instruction = "vssseg2e32.v,e8,mf8";
	    34'b0100111???????111?00010110?????001  :  Instruction = "vssseg2e64.v,e8,mf8";
	    34'b0100111???????000?00011010?????001  :  Instruction = "vssseg2e8.v,e8,mf4";
	    34'b0100111???????101?00011010?????001  :  Instruction = "vssseg2e16.v,e8,mf4";
	    34'b0100111???????110?00011010?????001  :  Instruction = "vssseg2e32.v,e8,mf4";
	    34'b0100111???????111?00011010?????001  :  Instruction = "vssseg2e64.v,e8,mf4";
	    34'b0100111???????000?00011110?????001  :  Instruction = "vssseg2e8.v,e8,mf2";
	    34'b0100111???????101?00011110?????001  :  Instruction = "vssseg2e16.v,e8,mf2";
	    34'b0100111???????110?00011110?????001  :  Instruction = "vssseg2e32.v,e8,mf2";
	    34'b0100111???????111?00011110?????001  :  Instruction = "vssseg2e64.v,e8,mf2";
	    34'b0100111???????000?00000010?????001  :  Instruction = "vssseg2e8.v,e8,m1";
	    34'b0100111???????101?00000010?????001  :  Instruction = "vssseg2e16.v,e8,m1";
	    34'b0100111???????110?00000010?????001  :  Instruction = "vssseg2e32.v,e8,m1";
	    34'b0100111???????000?00000110?????001  :  Instruction = "vssseg2e8.v,e8,m2";
	    34'b0100111???????101?00000110?????001  :  Instruction = "vssseg2e16.v,e8,m2";
	    34'b0100111???????000?00001010?????001  :  Instruction = "vssseg2e8.v,e8,m4";
	    34'b0100111???????000?000101?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e8,mf8";
	    34'b0100111???????101?000101?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e8,mf8";
	    34'b0100111???????110?000101?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e8,mf8";
	    34'b0100111???????111?000101?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e8,mf8";
	    34'b0100111???????000?000110?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e8,mf4";
	    34'b0100111???????101?000110?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e8,mf4";
	    34'b0100111???????110?000110?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e8,mf4";
	    34'b0100111???????111?000110?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e8,mf4";
	    34'b0100111???????000?000111?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e8,mf2";
	    34'b0100111???????101?000111?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e8,mf2";
	    34'b0100111???????110?000111?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e8,mf2";
	    34'b0100111???????111?000111?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e8,mf2";
	    34'b0100111???????000?000000?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e8,m1";
	    34'b0100111???????101?000000?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e8,m1";
	    34'b0100111???????110?000000?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e8,m1";
	    34'b0100111???????111?000000?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e8,m1";
	    34'b0100111???????000?000001?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e8,m2";
	    34'b0100111???????101?000001?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e8,m2";
	    34'b0100111???????110?000001?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e8,m2";
	    34'b0100111???????000?000010?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e8,m4";
	    34'b0100111???????101?000010?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e8,m4";
	    34'b0100111???????000?00010100?0000010  :  Instruction = "vsseg3e8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000010  :  Instruction = "vsseg3e16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000010  :  Instruction = "vsseg3e32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000010  :  Instruction = "vsseg3e64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000010  :  Instruction = "vsseg3e8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000010  :  Instruction = "vsseg3e16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000010  :  Instruction = "vsseg3e32[ff].v,e8,mf4";
	    34'b0100111???????111?00011000?0000010  :  Instruction = "vsseg3e64[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000010  :  Instruction = "vsseg3e8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000010  :  Instruction = "vsseg3e16[ff].v,e8,mf2";
	    34'b0100111???????110?00011100?0000010  :  Instruction = "vsseg3e32[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000010  :  Instruction = "vsseg3e8[ff].v,e8,m1";
	    34'b0100111???????101?00000000?0000010  :  Instruction = "vsseg3e16[ff].v,e8,m1";
	    34'b0100111???????000?00000100?0000010  :  Instruction = "vsseg3e8[ff].v,e8,m2";
	    34'b0100111???????000?00010110?????010  :  Instruction = "vssseg3e8.v,e8,mf8";
	    34'b0100111???????101?00010110?????010  :  Instruction = "vssseg3e16.v,e8,mf8";
	    34'b0100111???????110?00010110?????010  :  Instruction = "vssseg3e32.v,e8,mf8";
	    34'b0100111???????111?00010110?????010  :  Instruction = "vssseg3e64.v,e8,mf8";
	    34'b0100111???????000?00011010?????010  :  Instruction = "vssseg3e8.v,e8,mf4";
	    34'b0100111???????101?00011010?????010  :  Instruction = "vssseg3e16.v,e8,mf4";
	    34'b0100111???????110?00011010?????010  :  Instruction = "vssseg3e32.v,e8,mf4";
	    34'b0100111???????111?00011010?????010  :  Instruction = "vssseg3e64.v,e8,mf4";
	    34'b0100111???????000?00011110?????010  :  Instruction = "vssseg3e8.v,e8,mf2";
	    34'b0100111???????101?00011110?????010  :  Instruction = "vssseg3e16.v,e8,mf2";
	    34'b0100111???????110?00011110?????010  :  Instruction = "vssseg3e32.v,e8,mf2";
	    34'b0100111???????000?00000010?????010  :  Instruction = "vssseg3e8.v,e8,m1";
	    34'b0100111???????101?00000010?????010  :  Instruction = "vssseg3e16.v,e8,m1";
	    34'b0100111???????000?00000110?????010  :  Instruction = "vssseg3e8.v,e8,m2";
	    34'b0100111???????000?000101?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e8,mf8";
	    34'b0100111???????101?000101?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e8,mf8";
	    34'b0100111???????110?000101?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e8,mf8";
	    34'b0100111???????111?000101?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e8,mf8";
	    34'b0100111???????000?000110?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e8,mf4";
	    34'b0100111???????101?000110?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e8,mf4";
	    34'b0100111???????110?000110?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e8,mf4";
	    34'b0100111???????111?000110?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e8,mf4";
	    34'b0100111???????000?000111?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e8,mf2";
	    34'b0100111???????101?000111?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e8,mf2";
	    34'b0100111???????110?000111?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e8,mf2";
	    34'b0100111???????111?000111?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e8,mf2";
	    34'b0100111???????000?000000?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e8,m1";
	    34'b0100111???????101?000000?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e8,m1";
	    34'b0100111???????110?000000?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e8,m1";
	    34'b0100111???????111?000000?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e8,m1";
	    34'b0100111???????000?000001?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e8,m2";
	    34'b0100111???????101?000001?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e8,m2";
	    34'b0100111???????110?000001?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e8,m2";
	    34'b0100111???????000?00010100?0000011  :  Instruction = "vsseg4e8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000011  :  Instruction = "vsseg4e16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000011  :  Instruction = "vsseg4e32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000011  :  Instruction = "vsseg4e64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000011  :  Instruction = "vsseg4e8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000011  :  Instruction = "vsseg4e16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000011  :  Instruction = "vsseg4e32[ff].v,e8,mf4";
	    34'b0100111???????111?00011000?0000011  :  Instruction = "vsseg4e64[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000011  :  Instruction = "vsseg4e8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000011  :  Instruction = "vsseg4e16[ff].v,e8,mf2";
	    34'b0100111???????110?00011100?0000011  :  Instruction = "vsseg4e32[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000011  :  Instruction = "vsseg4e8[ff].v,e8,m1";
	    34'b0100111???????101?00000000?0000011  :  Instruction = "vsseg4e16[ff].v,e8,m1";
	    34'b0100111???????000?00000100?0000011  :  Instruction = "vsseg4e8[ff].v,e8,m2";
	    34'b0100111???????000?00010110?????011  :  Instruction = "vssseg4e8.v,e8,mf8";
	    34'b0100111???????101?00010110?????011  :  Instruction = "vssseg4e16.v,e8,mf8";
	    34'b0100111???????110?00010110?????011  :  Instruction = "vssseg4e32.v,e8,mf8";
	    34'b0100111???????111?00010110?????011  :  Instruction = "vssseg4e64.v,e8,mf8";
	    34'b0100111???????000?00011010?????011  :  Instruction = "vssseg4e8.v,e8,mf4";
	    34'b0100111???????101?00011010?????011  :  Instruction = "vssseg4e16.v,e8,mf4";
	    34'b0100111???????110?00011010?????011  :  Instruction = "vssseg4e32.v,e8,mf4";
	    34'b0100111???????111?00011010?????011  :  Instruction = "vssseg4e64.v,e8,mf4";
	    34'b0100111???????000?00011110?????011  :  Instruction = "vssseg4e8.v,e8,mf2";
	    34'b0100111???????101?00011110?????011  :  Instruction = "vssseg4e16.v,e8,mf2";
	    34'b0100111???????110?00011110?????011  :  Instruction = "vssseg4e32.v,e8,mf2";
	    34'b0100111???????000?00000010?????011  :  Instruction = "vssseg4e8.v,e8,m1";
	    34'b0100111???????101?00000010?????011  :  Instruction = "vssseg4e16.v,e8,m1";
	    34'b0100111???????000?00000110?????011  :  Instruction = "vssseg4e8.v,e8,m2";
	    34'b0100111???????000?000???0001000011  :  Instruction = "vs4r.v,e8";
	    34'b0100111???????000?000101?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e8,mf8";
	    34'b0100111???????101?000101?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e8,mf8";
	    34'b0100111???????110?000101?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e8,mf8";
	    34'b0100111???????111?000101?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e8,mf8";
	    34'b0100111???????000?000110?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e8,mf4";
	    34'b0100111???????101?000110?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e8,mf4";
	    34'b0100111???????110?000110?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e8,mf4";
	    34'b0100111???????111?000110?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e8,mf4";
	    34'b0100111???????000?000111?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e8,mf2";
	    34'b0100111???????101?000111?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e8,mf2";
	    34'b0100111???????110?000111?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e8,mf2";
	    34'b0100111???????111?000111?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e8,mf2";
	    34'b0100111???????000?000000?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e8,m1";
	    34'b0100111???????101?000000?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e8,m1";
	    34'b0100111???????110?000000?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e8,m1";
	    34'b0100111???????111?000000?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e8,m1";
	    34'b0100111???????000?000001?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e8,m2";
	    34'b0100111???????101?000001?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e8,m2";
	    34'b0100111???????110?000001?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e8,m2";
	    34'b0100111???????000?00010100?0000100  :  Instruction = "vsseg5e8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000100  :  Instruction = "vsseg5e16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000100  :  Instruction = "vsseg5e32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000100  :  Instruction = "vsseg5e64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000100  :  Instruction = "vsseg5e8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000100  :  Instruction = "vsseg5e16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000100  :  Instruction = "vsseg5e32[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000100  :  Instruction = "vsseg5e8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000100  :  Instruction = "vsseg5e16[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000100  :  Instruction = "vsseg5e8[ff].v,e8,m1";
	    34'b0100111???????000?00010110?????100  :  Instruction = "vssseg5e8.v,e8,mf8";
	    34'b0100111???????101?00010110?????100  :  Instruction = "vssseg5e16.v,e8,mf8";
	    34'b0100111???????110?00010110?????100  :  Instruction = "vssseg5e32.v,e8,mf8";
	    34'b0100111???????111?00010110?????100  :  Instruction = "vssseg5e64.v,e8,mf8";
	    34'b0100111???????000?00011010?????100  :  Instruction = "vssseg5e8.v,e8,mf4";
	    34'b0100111???????101?00011010?????100  :  Instruction = "vssseg5e16.v,e8,mf4";
	    34'b0100111???????110?00011010?????100  :  Instruction = "vssseg5e32.v,e8,mf4";
	    34'b0100111???????000?00011110?????100  :  Instruction = "vssseg5e8.v,e8,mf2";
	    34'b0100111???????101?00011110?????100  :  Instruction = "vssseg5e16.v,e8,mf2";
	    34'b0100111???????000?00000010?????100  :  Instruction = "vssseg5e8.v,e8,m1";
	    34'b0100111???????000?000101?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e8,mf8";
	    34'b0100111???????101?000101?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e8,mf8";
	    34'b0100111???????110?000101?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e8,mf8";
	    34'b0100111???????111?000101?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e8,mf8";
	    34'b0100111???????000?000110?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e8,mf4";
	    34'b0100111???????101?000110?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e8,mf4";
	    34'b0100111???????110?000110?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e8,mf4";
	    34'b0100111???????111?000110?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e8,mf4";
	    34'b0100111???????000?000111?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e8,mf2";
	    34'b0100111???????101?000111?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e8,mf2";
	    34'b0100111???????110?000111?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e8,mf2";
	    34'b0100111???????111?000111?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e8,mf2";
	    34'b0100111???????000?000000?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e8,m1";
	    34'b0100111???????101?000000?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e8,m1";
	    34'b0100111???????110?000000?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e8,m1";
	    34'b0100111???????111?000000?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e8,m1";
	    34'b0100111???????000?00010100?0000101  :  Instruction = "vsseg6e8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000101  :  Instruction = "vsseg6e16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000101  :  Instruction = "vsseg6e32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000101  :  Instruction = "vsseg6e64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000101  :  Instruction = "vsseg6e8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000101  :  Instruction = "vsseg6e16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000101  :  Instruction = "vsseg6e32[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000101  :  Instruction = "vsseg6e8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000101  :  Instruction = "vsseg6e16[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000101  :  Instruction = "vsseg6e8[ff].v,e8,m1";
	    34'b0100111???????000?00010110?????101  :  Instruction = "vssseg6e8.v,e8,mf8";
	    34'b0100111???????101?00010110?????101  :  Instruction = "vssseg6e16.v,e8,mf8";
	    34'b0100111???????110?00010110?????101  :  Instruction = "vssseg6e32.v,e8,mf8";
	    34'b0100111???????111?00010110?????101  :  Instruction = "vssseg6e64.v,e8,mf8";
	    34'b0100111???????000?00011010?????101  :  Instruction = "vssseg6e8.v,e8,mf4";
	    34'b0100111???????101?00011010?????101  :  Instruction = "vssseg6e16.v,e8,mf4";
	    34'b0100111???????110?00011010?????101  :  Instruction = "vssseg6e32.v,e8,mf4";
	    34'b0100111???????000?00011110?????101  :  Instruction = "vssseg6e8.v,e8,mf2";
	    34'b0100111???????101?00011110?????101  :  Instruction = "vssseg6e16.v,e8,mf2";
	    34'b0100111???????000?00000010?????101  :  Instruction = "vssseg6e8.v,e8,m1";
	    34'b0100111???????000?000101?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e8,mf8";
	    34'b0100111???????101?000101?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e8,mf8";
	    34'b0100111???????110?000101?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e8,mf8";
	    34'b0100111???????111?000101?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e8,mf8";
	    34'b0100111???????000?000110?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e8,mf4";
	    34'b0100111???????101?000110?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e8,mf4";
	    34'b0100111???????110?000110?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e8,mf4";
	    34'b0100111???????111?000110?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e8,mf4";
	    34'b0100111???????000?000111?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e8,mf2";
	    34'b0100111???????101?000111?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e8,mf2";
	    34'b0100111???????110?000111?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e8,mf2";
	    34'b0100111???????111?000111?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e8,mf2";
	    34'b0100111???????000?000000?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e8,m1";
	    34'b0100111???????101?000000?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e8,m1";
	    34'b0100111???????110?000000?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e8,m1";
	    34'b0100111???????111?000000?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e8,m1";
	    34'b0100111???????000?00010100?0000110  :  Instruction = "vsseg7e8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000110  :  Instruction = "vsseg7e16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000110  :  Instruction = "vsseg7e32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000110  :  Instruction = "vsseg7e64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000110  :  Instruction = "vsseg7e8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000110  :  Instruction = "vsseg7e16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000110  :  Instruction = "vsseg7e32[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000110  :  Instruction = "vsseg7e8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000110  :  Instruction = "vsseg7e16[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000110  :  Instruction = "vsseg7e8[ff].v,e8,m1";
	    34'b0100111???????000?00010110?????110  :  Instruction = "vssseg7e8.v,e8,mf8";
	    34'b0100111???????101?00010110?????110  :  Instruction = "vssseg7e16.v,e8,mf8";
	    34'b0100111???????110?00010110?????110  :  Instruction = "vssseg7e32.v,e8,mf8";
	    34'b0100111???????111?00010110?????110  :  Instruction = "vssseg7e64.v,e8,mf8";
	    34'b0100111???????000?00011010?????110  :  Instruction = "vssseg7e8.v,e8,mf4";
	    34'b0100111???????101?00011010?????110  :  Instruction = "vssseg7e16.v,e8,mf4";
	    34'b0100111???????110?00011010?????110  :  Instruction = "vssseg7e32.v,e8,mf4";
	    34'b0100111???????000?00011110?????110  :  Instruction = "vssseg7e8.v,e8,mf2";
	    34'b0100111???????101?00011110?????110  :  Instruction = "vssseg7e16.v,e8,mf2";
	    34'b0100111???????000?00000010?????110  :  Instruction = "vssseg7e8.v,e8,m1";
	    34'b0100111???????000?000101?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e8,mf8";
	    34'b0100111???????101?000101?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e8,mf8";
	    34'b0100111???????110?000101?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e8,mf8";
	    34'b0100111???????111?000101?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e8,mf8";
	    34'b0100111???????000?000110?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e8,mf4";
	    34'b0100111???????101?000110?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e8,mf4";
	    34'b0100111???????110?000110?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e8,mf4";
	    34'b0100111???????111?000110?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e8,mf4";
	    34'b0100111???????000?000111?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e8,mf2";
	    34'b0100111???????101?000111?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e8,mf2";
	    34'b0100111???????110?000111?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e8,mf2";
	    34'b0100111???????111?000111?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e8,mf2";
	    34'b0100111???????000?000000?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e8,m1";
	    34'b0100111???????101?000000?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e8,m1";
	    34'b0100111???????110?000000?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e8,m1";
	    34'b0100111???????111?000000?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e8,m1";
	    34'b0100111???????000?00010100?0000111  :  Instruction = "vsseg8e8[ff].v,e8,mf8";
	    34'b0100111???????101?00010100?0000111  :  Instruction = "vsseg8e16[ff].v,e8,mf8";
	    34'b0100111???????110?00010100?0000111  :  Instruction = "vsseg8e32[ff].v,e8,mf8";
	    34'b0100111???????111?00010100?0000111  :  Instruction = "vsseg8e64[ff].v,e8,mf8";
	    34'b0100111???????000?00011000?0000111  :  Instruction = "vsseg8e8[ff].v,e8,mf4";
	    34'b0100111???????101?00011000?0000111  :  Instruction = "vsseg8e16[ff].v,e8,mf4";
	    34'b0100111???????110?00011000?0000111  :  Instruction = "vsseg8e32[ff].v,e8,mf4";
	    34'b0100111???????000?00011100?0000111  :  Instruction = "vsseg8e8[ff].v,e8,mf2";
	    34'b0100111???????101?00011100?0000111  :  Instruction = "vsseg8e16[ff].v,e8,mf2";
	    34'b0100111???????000?00000000?0000111  :  Instruction = "vsseg8e8[ff].v,e8,m1";
	    34'b0100111???????000?000???0001000111  :  Instruction = "vs8r.v,e8";
	    34'b0100111???????000?00010110?????111  :  Instruction = "vssseg8e8.v,e8,mf8";
	    34'b0100111???????101?00010110?????111  :  Instruction = "vssseg8e16.v,e8,mf8";
	    34'b0100111???????110?00010110?????111  :  Instruction = "vssseg8e32.v,e8,mf8";
	    34'b0100111???????111?00010110?????111  :  Instruction = "vssseg8e64.v,e8,mf8";
	    34'b0100111???????000?00011010?????111  :  Instruction = "vssseg8e8.v,e8,mf4";
	    34'b0100111???????101?00011010?????111  :  Instruction = "vssseg8e16.v,e8,mf4";
	    34'b0100111???????110?00011010?????111  :  Instruction = "vssseg8e32.v,e8,mf4";
	    34'b0100111???????000?00011110?????111  :  Instruction = "vssseg8e8.v,e8,mf2";
	    34'b0100111???????101?00011110?????111  :  Instruction = "vssseg8e16.v,e8,mf2";
	    34'b0100111???????000?00000010?????111  :  Instruction = "vssseg8e8.v,e8,m1";
	    34'b0100111???????000?000101?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e8,mf8";
	    34'b0100111???????101?000101?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e8,mf8";
	    34'b0100111???????110?000101?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e8,mf8";
	    34'b0100111???????111?000101?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e8,mf8";
	    34'b0100111???????000?000110?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e8,mf4";
	    34'b0100111???????101?000110?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e8,mf4";
	    34'b0100111???????110?000110?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e8,mf4";
	    34'b0100111???????111?000110?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e8,mf4";
	    34'b0100111???????000?000111?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e8,mf2";
	    34'b0100111???????101?000111?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e8,mf2";
	    34'b0100111???????110?000111?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e8,mf2";
	    34'b0100111???????111?000111?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e8,mf2";
	    34'b0100111???????000?000000?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e8,m1";
	    34'b0100111???????101?000000?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e8,m1";
	    34'b0100111???????110?000000?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e8,m1";
	    34'b0100111???????111?000000?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e8,m1";
	    34'b0000111???????101?00110100?0000???  :  Instruction = "vle16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000???  :  Instruction = "vle32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000???  :  Instruction = "vle64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000???  :  Instruction = "vle8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000???  :  Instruction = "vle16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000???  :  Instruction = "vle32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000???  :  Instruction = "vle64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000???  :  Instruction = "vle8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000???  :  Instruction = "vle16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000???  :  Instruction = "vle32[ff].v,e16,mf2";
	    34'b0000111???????111?00111100?0000???  :  Instruction = "vle64[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000???  :  Instruction = "vle8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000???  :  Instruction = "vle16[ff].v,e16,m1";
	    34'b0000111???????110?00100000?0000???  :  Instruction = "vle32[ff].v,e16,m1";
	    34'b0000111???????111?00100000?0000???  :  Instruction = "vle64[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000???  :  Instruction = "vle8[ff].v,e16,m2";
	    34'b0000111???????101?00100100?0000???  :  Instruction = "vle16[ff].v,e16,m2";
	    34'b0000111???????110?00100100?0000???  :  Instruction = "vle32[ff].v,e16,m2";
	    34'b0000111???????111?00100100?0000???  :  Instruction = "vle64[ff].v,e16,m2";
	    34'b0000111???????000?00101000?0000???  :  Instruction = "vle8[ff].v,e16,m4";
	    34'b0000111???????101?00101000?0000???  :  Instruction = "vle16[ff].v,e16,m4";
	    34'b0000111???????110?00101000?0000???  :  Instruction = "vle32[ff].v,e16,m4";
	    34'b0000111???????000?00101100?0000???  :  Instruction = "vle8[ff].v,e16,m8";
	    34'b0000111???????101?00101100?0000???  :  Instruction = "vle16[ff].v,e16,m8";
	    34'b0000111???????000?001???0001000000  :  Instruction = "vl1re8.v,e16";
	    34'b0000111???????101?001???0001000000  :  Instruction = "vl1re16.v,e16";
	    34'b0000111???????110?001???0001000000  :  Instruction = "vl1re32.v,e16";
	    34'b0000111???????111?001???0001000000  :  Instruction = "vl1re64.v,e16";
	    34'b0000111???????101?00110110????????  :  Instruction = "vlse16.v,e16,mf8";
	    34'b0000111???????110?00110110????????  :  Instruction = "vlse32.v,e16,mf8";
	    34'b0000111???????111?00110110????????  :  Instruction = "vlse64.v,e16,mf8";
	    34'b0000111???????000?00111010????????  :  Instruction = "vlse8.v,e16,mf4";
	    34'b0000111???????101?00111010????????  :  Instruction = "vlse16.v,e16,mf4";
	    34'b0000111???????110?00111010????????  :  Instruction = "vlse32.v,e16,mf4";
	    34'b0000111???????111?00111010????????  :  Instruction = "vlse64.v,e16,mf4";
	    34'b0000111???????000?00111110????????  :  Instruction = "vlse8.v,e16,mf2";
	    34'b0000111???????101?00111110????????  :  Instruction = "vlse16.v,e16,mf2";
	    34'b0000111???????110?00111110????????  :  Instruction = "vlse32.v,e16,mf2";
	    34'b0000111???????111?00111110????????  :  Instruction = "vlse64.v,e16,mf2";
	    34'b0000111???????000?00100010????????  :  Instruction = "vlse8.v,e16,m1";
	    34'b0000111???????101?00100010????????  :  Instruction = "vlse16.v,e16,m1";
	    34'b0000111???????110?00100010????????  :  Instruction = "vlse32.v,e16,m1";
	    34'b0000111???????111?00100010????????  :  Instruction = "vlse64.v,e16,m1";
	    34'b0000111???????000?00100110????????  :  Instruction = "vlse8.v,e16,m2";
	    34'b0000111???????101?00100110????????  :  Instruction = "vlse16.v,e16,m2";
	    34'b0000111???????110?00100110????????  :  Instruction = "vlse32.v,e16,m2";
	    34'b0000111???????111?00100110????????  :  Instruction = "vlse64.v,e16,m2";
	    34'b0000111???????000?00101010????????  :  Instruction = "vlse8.v,e16,m4";
	    34'b0000111???????101?00101010????????  :  Instruction = "vlse16.v,e16,m4";
	    34'b0000111???????110?00101010????????  :  Instruction = "vlse32.v,e16,m4";
	    34'b0000111???????000?00101110????????  :  Instruction = "vlse8.v,e16,m8";
	    34'b0000111???????101?00101110????????  :  Instruction = "vlse16.v,e16,m8";
	    34'b0000111???????101?001101?1????????  :  Instruction = "vl[uo]xei16.v,e16,mf8";
	    34'b0000111???????110?001101?1????????  :  Instruction = "vl[uo]xei32.v,e16,mf8";
	    34'b0000111???????111?001101?1????????  :  Instruction = "vl[uo]xei64.v,e16,mf8";
	    34'b0000111???????000?001110?1????????  :  Instruction = "vl[uo]xei8.v,e16,mf4";
	    34'b0000111???????101?001110?1????????  :  Instruction = "vl[uo]xei16.v,e16,mf4";
	    34'b0000111???????110?001110?1????????  :  Instruction = "vl[uo]xei32.v,e16,mf4";
	    34'b0000111???????111?001110?1????????  :  Instruction = "vl[uo]xei64.v,e16,mf4";
	    34'b0000111???????000?001111?1????????  :  Instruction = "vl[uo]xei8.v,e16,mf2";
	    34'b0000111???????101?001111?1????????  :  Instruction = "vl[uo]xei16.v,e16,mf2";
	    34'b0000111???????110?001111?1????????  :  Instruction = "vl[uo]xei32.v,e16,mf2";
	    34'b0000111???????111?001111?1????????  :  Instruction = "vl[uo]xei64.v,e16,mf2";
	    34'b0000111???????000?001000?1????????  :  Instruction = "vl[uo]xei8.v,e16,m1";
	    34'b0000111???????101?001000?1????????  :  Instruction = "vl[uo]xei16.v,e16,m1";
	    34'b0000111???????110?001000?1????????  :  Instruction = "vl[uo]xei32.v,e16,m1";
	    34'b0000111???????111?001000?1????????  :  Instruction = "vl[uo]xei64.v,e16,m1";
	    34'b0000111???????000?001001?1????????  :  Instruction = "vl[uo]xei8.v,e16,m2";
	    34'b0000111???????101?001001?1????????  :  Instruction = "vl[uo]xei16.v,e16,m2";
	    34'b0000111???????110?001001?1????????  :  Instruction = "vl[uo]xei32.v,e16,m2";
	    34'b0000111???????111?001001?1????????  :  Instruction = "vl[uo]xei64.v,e16,m2";
	    34'b0000111???????000?001010?1????????  :  Instruction = "vl[uo]xei8.v,e16,m4";
	    34'b0000111???????101?001010?1????????  :  Instruction = "vl[uo]xei16.v,e16,m4";
	    34'b0000111???????110?001010?1????????  :  Instruction = "vl[uo]xei32.v,e16,m4";
	    34'b0000111???????000?001011?1????????  :  Instruction = "vl[uo]xei8.v,e16,m8";
	    34'b0000111???????101?001011?1????????  :  Instruction = "vl[uo]xei16.v,e16,m8";
	    34'b0000111???????101?00110100?0000001  :  Instruction = "vlseg2e16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000001  :  Instruction = "vlseg2e32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000001  :  Instruction = "vlseg2e64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000001  :  Instruction = "vlseg2e8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000001  :  Instruction = "vlseg2e16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000001  :  Instruction = "vlseg2e32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000001  :  Instruction = "vlseg2e64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000001  :  Instruction = "vlseg2e8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000001  :  Instruction = "vlseg2e16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000001  :  Instruction = "vlseg2e32[ff].v,e16,mf2";
	    34'b0000111???????111?00111100?0000001  :  Instruction = "vlseg2e64[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000001  :  Instruction = "vlseg2e8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000001  :  Instruction = "vlseg2e16[ff].v,e16,m1";
	    34'b0000111???????110?00100000?0000001  :  Instruction = "vlseg2e32[ff].v,e16,m1";
	    34'b0000111???????111?00100000?0000001  :  Instruction = "vlseg2e64[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000001  :  Instruction = "vlseg2e8[ff].v,e16,m2";
	    34'b0000111???????101?00100100?0000001  :  Instruction = "vlseg2e16[ff].v,e16,m2";
	    34'b0000111???????110?00100100?0000001  :  Instruction = "vlseg2e32[ff].v,e16,m2";
	    34'b0000111???????000?00101000?0000001  :  Instruction = "vlseg2e8[ff].v,e16,m4";
	    34'b0000111???????101?00101000?0000001  :  Instruction = "vlseg2e16[ff].v,e16,m4";
	    34'b0000111???????000?00101100?0000001  :  Instruction = "vlseg2e8[ff].v,e16,m8";
	    34'b0000111???????111?00101100?0000001  :  Instruction = "vlseg2e64[ff].v,e16,m8";
	    34'b0000111???????000?001???0001000001  :  Instruction = "vl2re8.v,e16";
	    34'b0000111???????101?001???0001000001  :  Instruction = "vl2re16.v,e16";
	    34'b0000111???????110?001???0001000001  :  Instruction = "vl2re32.v,e16";
	    34'b0000111???????111?001???0001000001  :  Instruction = "vl2re64.v,e16";
	    34'b0000111???????101?00110110?????001  :  Instruction = "vlsseg2e16.v,e16,mf8";
	    34'b0000111???????110?00110110?????001  :  Instruction = "vlsseg2e32.v,e16,mf8";
	    34'b0000111???????111?00110110?????001  :  Instruction = "vlsseg2e64.v,e16,mf8";
	    34'b0000111???????000?00111010?????001  :  Instruction = "vlsseg2e8.v,e16,mf4";
	    34'b0000111???????101?00111010?????001  :  Instruction = "vlsseg2e16.v,e16,mf4";
	    34'b0000111???????110?00111010?????001  :  Instruction = "vlsseg2e32.v,e16,mf4";
	    34'b0000111???????111?00111010?????001  :  Instruction = "vlsseg2e64.v,e16,mf4";
	    34'b0000111???????000?00111110?????001  :  Instruction = "vlsseg2e8.v,e16,mf2";
	    34'b0000111???????101?00111110?????001  :  Instruction = "vlsseg2e16.v,e16,mf2";
	    34'b0000111???????110?00111110?????001  :  Instruction = "vlsseg2e32.v,e16,mf2";
	    34'b0000111???????111?00111110?????001  :  Instruction = "vlsseg2e64.v,e16,mf2";
	    34'b0000111???????000?00100010?????001  :  Instruction = "vlsseg2e8.v,e16,m1";
	    34'b0000111???????101?00100010?????001  :  Instruction = "vlsseg2e16.v,e16,m1";
	    34'b0000111???????110?00100010?????001  :  Instruction = "vlsseg2e32.v,e16,m1";
	    34'b0000111???????111?00100010?????001  :  Instruction = "vlsseg2e64.v,e16,m1";
	    34'b0000111???????000?00100110?????001  :  Instruction = "vlsseg2e8.v,e16,m2";
	    34'b0000111???????101?00100110?????001  :  Instruction = "vlsseg2e16.v,e16,m2";
	    34'b0000111???????110?00100110?????001  :  Instruction = "vlsseg2e32.v,e16,m2";
	    34'b0000111???????000?00101010?????001  :  Instruction = "vlsseg2e8.v,e16,m4";
	    34'b0000111???????101?00101010?????001  :  Instruction = "vlsseg2e16.v,e16,m4";
	    34'b0000111???????000?00101110?????001  :  Instruction = "vlsseg2e8.v,e16,m8";
	    34'b0000111???????101?001101?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e16,mf8";
	    34'b0000111???????110?001101?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e16,mf8";
	    34'b0000111???????111?001101?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e16,mf8";
	    34'b0000111???????000?001110?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e16,mf4";
	    34'b0000111???????101?001110?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e16,mf4";
	    34'b0000111???????110?001110?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e16,mf4";
	    34'b0000111???????111?001110?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e16,mf4";
	    34'b0000111???????000?001111?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e16,mf2";
	    34'b0000111???????101?001111?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e16,mf2";
	    34'b0000111???????110?001111?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e16,mf2";
	    34'b0000111???????111?001111?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e16,mf2";
	    34'b0000111???????000?001000?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e16,m1";
	    34'b0000111???????101?001000?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e16,m1";
	    34'b0000111???????110?001000?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e16,m1";
	    34'b0000111???????111?001000?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e16,m1";
	    34'b0000111???????000?001001?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e16,m2";
	    34'b0000111???????101?001001?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e16,m2";
	    34'b0000111???????110?001001?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e16,m2";
	    34'b0000111???????111?001001?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e16,m2";
	    34'b0000111???????000?001010?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e16,m4";
	    34'b0000111???????101?001010?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e16,m4";
	    34'b0000111???????110?001010?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e16,m4";
	    34'b0000111???????101?00110100?0000010  :  Instruction = "vlseg3e16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000010  :  Instruction = "vlseg3e32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000010  :  Instruction = "vlseg3e64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000010  :  Instruction = "vlseg3e8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000010  :  Instruction = "vlseg3e16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000010  :  Instruction = "vlseg3e32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000010  :  Instruction = "vlseg3e64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000010  :  Instruction = "vlseg3e8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000010  :  Instruction = "vlseg3e16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000010  :  Instruction = "vlseg3e32[ff].v,e16,mf2";
	    34'b0000111???????111?00111100?0000010  :  Instruction = "vlseg3e64[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000010  :  Instruction = "vlseg3e8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000010  :  Instruction = "vlseg3e16[ff].v,e16,m1";
	    34'b0000111???????110?00100000?0000010  :  Instruction = "vlseg3e32[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000010  :  Instruction = "vlseg3e8[ff].v,e16,m2";
	    34'b0000111???????101?00100100?0000010  :  Instruction = "vlseg3e16[ff].v,e16,m2";
	    34'b0000111???????000?00101000?0000010  :  Instruction = "vlseg3e8[ff].v,e16,m4";
	    34'b0000111???????101?00110110?????010  :  Instruction = "vlsseg3e16.v,e16,mf8";
	    34'b0000111???????110?00110110?????010  :  Instruction = "vlsseg3e32.v,e16,mf8";
	    34'b0000111???????111?00110110?????010  :  Instruction = "vlsseg3e64.v,e16,mf8";
	    34'b0000111???????000?00111010?????010  :  Instruction = "vlsseg3e8.v,e16,mf4";
	    34'b0000111???????101?00111010?????010  :  Instruction = "vlsseg3e16.v,e16,mf4";
	    34'b0000111???????110?00111010?????010  :  Instruction = "vlsseg3e32.v,e16,mf4";
	    34'b0000111???????111?00111010?????010  :  Instruction = "vlsseg3e64.v,e16,mf4";
	    34'b0000111???????000?00111110?????010  :  Instruction = "vlsseg3e8.v,e16,mf2";
	    34'b0000111???????101?00111110?????010  :  Instruction = "vlsseg3e16.v,e16,mf2";
	    34'b0000111???????110?00111110?????010  :  Instruction = "vlsseg3e32.v,e16,mf2";
	    34'b0000111???????111?00111110?????010  :  Instruction = "vlsseg3e64.v,e16,mf2";
	    34'b0000111???????000?00100010?????010  :  Instruction = "vlsseg3e8.v,e16,m1";
	    34'b0000111???????101?00100010?????010  :  Instruction = "vlsseg3e16.v,e16,m1";
	    34'b0000111???????110?00100010?????010  :  Instruction = "vlsseg3e32.v,e16,m1";
	    34'b0000111???????000?00100110?????010  :  Instruction = "vlsseg3e8.v,e16,m2";
	    34'b0000111???????101?00100110?????010  :  Instruction = "vlsseg3e16.v,e16,m2";
	    34'b0000111???????000?00101010?????010  :  Instruction = "vlsseg3e8.v,e16,m4";
	    34'b0000111???????101?001101?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e16,mf8";
	    34'b0000111???????110?001101?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e16,mf8";
	    34'b0000111???????111?001101?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e16,mf8";
	    34'b0000111???????000?001110?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e16,mf4";
	    34'b0000111???????101?001110?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e16,mf4";
	    34'b0000111???????110?001110?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e16,mf4";
	    34'b0000111???????111?001110?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e16,mf4";
	    34'b0000111???????000?001111?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e16,mf2";
	    34'b0000111???????101?001111?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e16,mf2";
	    34'b0000111???????110?001111?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e16,mf2";
	    34'b0000111???????111?001111?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e16,mf2";
	    34'b0000111???????000?001000?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e16,m1";
	    34'b0000111???????101?001000?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e16,m1";
	    34'b0000111???????110?001000?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e16,m1";
	    34'b0000111???????111?001000?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e16,m1";
	    34'b0000111???????000?001001?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e16,m2";
	    34'b0000111???????101?001001?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e16,m2";
	    34'b0000111???????110?001001?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e16,m2";
	    34'b0000111???????111?001001?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e16,m2";
	    34'b0000111???????101?00110100?0000011  :  Instruction = "vlseg4e16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000011  :  Instruction = "vlseg4e32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000011  :  Instruction = "vlseg4e64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000011  :  Instruction = "vlseg4e8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000011  :  Instruction = "vlseg4e16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000011  :  Instruction = "vlseg4e32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000011  :  Instruction = "vlseg4e64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000011  :  Instruction = "vlseg4e8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000011  :  Instruction = "vlseg4e16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000011  :  Instruction = "vlseg4e32[ff].v,e16,mf2";
	    34'b0000111???????111?00111100?0000011  :  Instruction = "vlseg4e64[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000011  :  Instruction = "vlseg4e8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000011  :  Instruction = "vlseg4e16[ff].v,e16,m1";
	    34'b0000111???????110?00100000?0000011  :  Instruction = "vlseg4e32[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000011  :  Instruction = "vlseg4e8[ff].v,e16,m2";
	    34'b0000111???????101?00100100?0000011  :  Instruction = "vlseg4e16[ff].v,e16,m2";
	    34'b0000111???????000?00101000?0000011  :  Instruction = "vlseg4e8[ff].v,e16,m4";
	    34'b0000111???????101?00110110?????011  :  Instruction = "vlsseg4e16.v,e16,mf8";
	    34'b0000111???????110?00110110?????011  :  Instruction = "vlsseg4e32.v,e16,mf8";
	    34'b0000111???????111?00110110?????011  :  Instruction = "vlsseg4e64.v,e16,mf8";
	    34'b0000111???????000?00111010?????011  :  Instruction = "vlsseg4e8.v,e16,mf4";
	    34'b0000111???????101?00111010?????011  :  Instruction = "vlsseg4e16.v,e16,mf4";
	    34'b0000111???????110?00111010?????011  :  Instruction = "vlsseg4e32.v,e16,mf4";
	    34'b0000111???????111?00111010?????011  :  Instruction = "vlsseg4e64.v,e16,mf4";
	    34'b0000111???????000?00111110?????011  :  Instruction = "vlsseg4e8.v,e16,mf2";
	    34'b0000111???????101?00111110?????011  :  Instruction = "vlsseg4e16.v,e16,mf2";
	    34'b0000111???????110?00111110?????011  :  Instruction = "vlsseg4e32.v,e16,mf2";
	    34'b0000111???????111?00111110?????011  :  Instruction = "vlsseg4e64.v,e16,mf2";
	    34'b0000111???????000?00100010?????011  :  Instruction = "vlsseg4e8.v,e16,m1";
	    34'b0000111???????101?00100010?????011  :  Instruction = "vlsseg4e16.v,e16,m1";
	    34'b0000111???????110?00100010?????011  :  Instruction = "vlsseg4e32.v,e16,m1";
	    34'b0000111???????000?00100110?????011  :  Instruction = "vlsseg4e8.v,e16,m2";
	    34'b0000111???????101?00100110?????011  :  Instruction = "vlsseg4e16.v,e16,m2";
	    34'b0000111???????000?00101010?????011  :  Instruction = "vlsseg4e8.v,e16,m4";
	    34'b0000111???????000?001???0001000011  :  Instruction = "vl4re8.v,e16";
	    34'b0000111???????101?001???0001000011  :  Instruction = "vl4re16.v,e16";
	    34'b0000111???????110?001???0001000011  :  Instruction = "vl4re32.v,e16";
	    34'b0000111???????111?001???0001000011  :  Instruction = "vl4re64.v,e16";
	    34'b0000111???????101?001101?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e16,mf8";
	    34'b0000111???????110?001101?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e16,mf8";
	    34'b0000111???????111?001101?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e16,mf8";
	    34'b0000111???????000?001110?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e16,mf4";
	    34'b0000111???????101?001110?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e16,mf4";
	    34'b0000111???????110?001110?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e16,mf4";
	    34'b0000111???????111?001110?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e16,mf4";
	    34'b0000111???????000?001111?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e16,mf2";
	    34'b0000111???????101?001111?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e16,mf2";
	    34'b0000111???????110?001111?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e16,mf2";
	    34'b0000111???????111?001111?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e16,mf2";
	    34'b0000111???????000?001000?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e16,m1";
	    34'b0000111???????101?001000?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e16,m1";
	    34'b0000111???????110?001000?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e16,m1";
	    34'b0000111???????111?001000?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e16,m1";
	    34'b0000111???????000?001001?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e16,m2";
	    34'b0000111???????101?001001?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e16,m2";
	    34'b0000111???????110?001001?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e16,m2";
	    34'b0000111???????111?001001?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e16,m2";
	    34'b0000111???????101?00110100?0000100  :  Instruction = "vlseg5e16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000100  :  Instruction = "vlseg5e32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000100  :  Instruction = "vlseg5e64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000100  :  Instruction = "vlseg5e8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000100  :  Instruction = "vlseg5e16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000100  :  Instruction = "vlseg5e32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000100  :  Instruction = "vlseg5e64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000100  :  Instruction = "vlseg5e8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000100  :  Instruction = "vlseg5e16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000100  :  Instruction = "vlseg5e32[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000100  :  Instruction = "vlseg5e8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000100  :  Instruction = "vlseg5e16[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000100  :  Instruction = "vlseg5e8[ff].v,e16,m2";
	    34'b0000111???????101?00110110?????100  :  Instruction = "vlsseg5e16.v,e16,mf8";
	    34'b0000111???????110?00110110?????100  :  Instruction = "vlsseg5e32.v,e16,mf8";
	    34'b0000111???????111?00110110?????100  :  Instruction = "vlsseg5e64.v,e16,mf8";
	    34'b0000111???????000?00111010?????100  :  Instruction = "vlsseg5e8.v,e16,mf4";
	    34'b0000111???????101?00111010?????100  :  Instruction = "vlsseg5e16.v,e16,mf4";
	    34'b0000111???????110?00111010?????100  :  Instruction = "vlsseg5e32.v,e16,mf4";
	    34'b0000111???????111?00111010?????100  :  Instruction = "vlsseg5e64.v,e16,mf4";
	    34'b0000111???????000?00111110?????100  :  Instruction = "vlsseg5e8.v,e16,mf2";
	    34'b0000111???????101?00111110?????100  :  Instruction = "vlsseg5e16.v,e16,mf2";
	    34'b0000111???????110?00111110?????100  :  Instruction = "vlsseg5e32.v,e16,mf2";
	    34'b0000111???????000?00100010?????100  :  Instruction = "vlsseg5e8.v,e16,m1";
	    34'b0000111???????101?00100010?????100  :  Instruction = "vlsseg5e16.v,e16,m1";
	    34'b0000111???????000?00100110?????100  :  Instruction = "vlsseg5e8.v,e16,m2";
	    34'b0000111???????101?001101?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e16,mf8";
	    34'b0000111???????110?001101?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e16,mf8";
	    34'b0000111???????111?001101?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e16,mf8";
	    34'b0000111???????000?001110?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e16,mf4";
	    34'b0000111???????101?001110?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e16,mf4";
	    34'b0000111???????110?001110?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e16,mf4";
	    34'b0000111???????111?001110?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e16,mf4";
	    34'b0000111???????000?001111?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e16,mf2";
	    34'b0000111???????101?001111?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e16,mf2";
	    34'b0000111???????110?001111?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e16,mf2";
	    34'b0000111???????111?001111?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e16,mf2";
	    34'b0000111???????000?001000?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e16,m1";
	    34'b0000111???????101?001000?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e16,m1";
	    34'b0000111???????110?001000?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e16,m1";
	    34'b0000111???????111?001000?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e16,m1";
	    34'b0000111???????101?00110100?0000101  :  Instruction = "vlseg6e16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000101  :  Instruction = "vlseg6e32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000101  :  Instruction = "vlseg6e64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000101  :  Instruction = "vlseg6e8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000101  :  Instruction = "vlseg6e16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000101  :  Instruction = "vlseg6e32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000101  :  Instruction = "vlseg6e64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000101  :  Instruction = "vlseg6e8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000101  :  Instruction = "vlseg6e16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000101  :  Instruction = "vlseg6e32[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000101  :  Instruction = "vlseg6e8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000101  :  Instruction = "vlseg6e16[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000101  :  Instruction = "vlseg6e8[ff].v,e16,m2";
	    34'b0000111???????101?00110110?????101  :  Instruction = "vlsseg6e16.v,e16,mf8";
	    34'b0000111???????110?00110110?????101  :  Instruction = "vlsseg6e32.v,e16,mf8";
	    34'b0000111???????111?00110110?????101  :  Instruction = "vlsseg6e64.v,e16,mf8";
	    34'b0000111???????000?00111010?????101  :  Instruction = "vlsseg6e8.v,e16,mf4";
	    34'b0000111???????101?00111010?????101  :  Instruction = "vlsseg6e16.v,e16,mf4";
	    34'b0000111???????110?00111010?????101  :  Instruction = "vlsseg6e32.v,e16,mf4";
	    34'b0000111???????111?00111010?????101  :  Instruction = "vlsseg6e64.v,e16,mf4";
	    34'b0000111???????000?00111110?????101  :  Instruction = "vlsseg6e8.v,e16,mf2";
	    34'b0000111???????101?00111110?????101  :  Instruction = "vlsseg6e16.v,e16,mf2";
	    34'b0000111???????110?00111110?????101  :  Instruction = "vlsseg6e32.v,e16,mf2";
	    34'b0000111???????000?00100010?????101  :  Instruction = "vlsseg6e8.v,e16,m1";
	    34'b0000111???????101?00100010?????101  :  Instruction = "vlsseg6e16.v,e16,m1";
	    34'b0000111???????000?00100110?????101  :  Instruction = "vlsseg6e8.v,e16,m2";
	    34'b0000111???????101?001101?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e16,mf8";
	    34'b0000111???????110?001101?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e16,mf8";
	    34'b0000111???????111?001101?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e16,mf8";
	    34'b0000111???????000?001110?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e16,mf4";
	    34'b0000111???????101?001110?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e16,mf4";
	    34'b0000111???????110?001110?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e16,mf4";
	    34'b0000111???????111?001110?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e16,mf4";
	    34'b0000111???????000?001111?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e16,mf2";
	    34'b0000111???????101?001111?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e16,mf2";
	    34'b0000111???????110?001111?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e16,mf2";
	    34'b0000111???????111?001111?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e16,mf2";
	    34'b0000111???????000?001000?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e16,m1";
	    34'b0000111???????101?001000?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e16,m1";
	    34'b0000111???????110?001000?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e16,m1";
	    34'b0000111???????111?001000?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e16,m1";
	    34'b0000111???????101?00110100?0000110  :  Instruction = "vlseg7e16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000110  :  Instruction = "vlseg7e32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000110  :  Instruction = "vlseg7e64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000110  :  Instruction = "vlseg7e8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000110  :  Instruction = "vlseg7e16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000110  :  Instruction = "vlseg7e32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000110  :  Instruction = "vlseg7e64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000110  :  Instruction = "vlseg7e8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000110  :  Instruction = "vlseg7e16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000110  :  Instruction = "vlseg7e32[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000110  :  Instruction = "vlseg7e8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000110  :  Instruction = "vlseg7e16[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000110  :  Instruction = "vlseg7e8[ff].v,e16,m2";
	    34'b0000111???????101?00110110?????110  :  Instruction = "vlsseg7e16.v,e16,mf8";
	    34'b0000111???????110?00110110?????110  :  Instruction = "vlsseg7e32.v,e16,mf8";
	    34'b0000111???????111?00110110?????110  :  Instruction = "vlsseg7e64.v,e16,mf8";
	    34'b0000111???????000?00111010?????110  :  Instruction = "vlsseg7e8.v,e16,mf4";
	    34'b0000111???????101?00111010?????110  :  Instruction = "vlsseg7e16.v,e16,mf4";
	    34'b0000111???????110?00111010?????110  :  Instruction = "vlsseg7e32.v,e16,mf4";
	    34'b0000111???????111?00111010?????110  :  Instruction = "vlsseg7e64.v,e16,mf4";
	    34'b0000111???????000?00111110?????110  :  Instruction = "vlsseg7e8.v,e16,mf2";
	    34'b0000111???????101?00111110?????110  :  Instruction = "vlsseg7e16.v,e16,mf2";
	    34'b0000111???????110?00111110?????110  :  Instruction = "vlsseg7e32.v,e16,mf2";
	    34'b0000111???????111?00111110?????110  :  Instruction = "vlsseg7e64.v,e16,mf2";
	    34'b0000111???????000?00100010?????110  :  Instruction = "vlsseg7e8.v,e16,m1";
	    34'b0000111???????101?00100010?????110  :  Instruction = "vlsseg7e16.v,e16,m1";
	    34'b0000111???????000?00100110?????110  :  Instruction = "vlsseg7e8.v,e16,m2";
	    34'b0000111???????101?001101?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e16,mf8";
	    34'b0000111???????110?001101?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e16,mf8";
	    34'b0000111???????111?001101?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e16,mf8";
	    34'b0000111???????000?001110?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e16,mf4";
	    34'b0000111???????101?001110?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e16,mf4";
	    34'b0000111???????110?001110?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e16,mf4";
	    34'b0000111???????111?001110?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e16,mf4";
	    34'b0000111???????000?001111?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e16,mf2";
	    34'b0000111???????101?001111?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e16,mf2";
	    34'b0000111???????110?001111?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e16,mf2";
	    34'b0000111???????111?001111?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e16,mf2";
	    34'b0000111???????000?001000?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e16,m1";
	    34'b0000111???????101?001000?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e16,m1";
	    34'b0000111???????110?001000?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e16,m1";
	    34'b0000111???????111?001000?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e16,m1";
	    34'b0000111???????101?00110100?0000111  :  Instruction = "vlseg8e16[ff].v,e16,mf8";
	    34'b0000111???????110?00110100?0000111  :  Instruction = "vlseg8e32[ff].v,e16,mf8";
	    34'b0000111???????111?00110100?0000111  :  Instruction = "vlseg8e64[ff].v,e16,mf8";
	    34'b0000111???????000?00111000?0000111  :  Instruction = "vlseg8e8[ff].v,e16,mf4";
	    34'b0000111???????101?00111000?0000111  :  Instruction = "vlseg8e16[ff].v,e16,mf4";
	    34'b0000111???????110?00111000?0000111  :  Instruction = "vlseg8e32[ff].v,e16,mf4";
	    34'b0000111???????111?00111000?0000111  :  Instruction = "vlseg8e64[ff].v,e16,mf4";
	    34'b0000111???????000?00111100?0000111  :  Instruction = "vlseg8e8[ff].v,e16,mf2";
	    34'b0000111???????101?00111100?0000111  :  Instruction = "vlseg8e16[ff].v,e16,mf2";
	    34'b0000111???????110?00111100?0000111  :  Instruction = "vlseg8e32[ff].v,e16,mf2";
	    34'b0000111???????000?00100000?0000111  :  Instruction = "vlseg8e8[ff].v,e16,m1";
	    34'b0000111???????101?00100000?0000111  :  Instruction = "vlseg8e16[ff].v,e16,m1";
	    34'b0000111???????000?00100100?0000111  :  Instruction = "vlseg8e8[ff].v,e16,m2";
	    34'b0000111???????000?001???0001000111  :  Instruction = "vl8re8.v,e16";
	    34'b0000111???????101?001???0001000111  :  Instruction = "vl8re16.v,e16";
	    34'b0000111???????110?001???0001000111  :  Instruction = "vl8re32.v,e16";
	    34'b0000111???????111?001???0001000111  :  Instruction = "vl8re64.v,e16";
	    34'b0000111???????101?00110110?????111  :  Instruction = "vlsseg8e16.v,e16,mf8";
	    34'b0000111???????110?00110110?????111  :  Instruction = "vlsseg8e32.v,e16,mf8";
	    34'b0000111???????111?00110110?????111  :  Instruction = "vlsseg8e64.v,e16,mf8";
	    34'b0000111???????000?00111010?????111  :  Instruction = "vlsseg8e8.v,e16,mf4";
	    34'b0000111???????101?00111010?????111  :  Instruction = "vlsseg8e16.v,e16,mf4";
	    34'b0000111???????110?00111010?????111  :  Instruction = "vlsseg8e32.v,e16,mf4";
	    34'b0000111???????111?00111010?????111  :  Instruction = "vlsseg8e64.v,e16,mf4";
	    34'b0000111???????000?00111110?????111  :  Instruction = "vlsseg8e8.v,e16,mf2";
	    34'b0000111???????101?00111110?????111  :  Instruction = "vlsseg8e16.v,e16,mf2";
	    34'b0000111???????110?00111110?????111  :  Instruction = "vlsseg8e32.v,e16,mf2";
	    34'b0000111???????000?00100010?????111  :  Instruction = "vlsseg8e8.v,e16,m1";
	    34'b0000111???????101?00100010?????111  :  Instruction = "vlsseg8e16.v,e16,m1";
	    34'b0000111???????000?00100110?????111  :  Instruction = "vlsseg8e8.v,e16,m2";
	    34'b0000111???????101?001101?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e16,mf8";
	    34'b0000111???????110?001101?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e16,mf8";
	    34'b0000111???????111?001101?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e16,mf8";
	    34'b0000111???????000?001110?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e16,mf4";
	    34'b0000111???????101?001110?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e16,mf4";
	    34'b0000111???????110?001110?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e16,mf4";
	    34'b0000111???????111?001110?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e16,mf4";
	    34'b0000111???????000?001111?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e16,mf2";
	    34'b0000111???????101?001111?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e16,mf2";
	    34'b0000111???????110?001111?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e16,mf2";
	    34'b0000111???????111?001111?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e16,mf2";
	    34'b0000111???????000?001000?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e16,m1";
	    34'b0000111???????101?001000?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e16,m1";
	    34'b0000111???????110?001000?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e16,m1";
	    34'b0000111???????111?001000?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e16,m1";
	    34'b0100111???????101?00110100?0000???  :  Instruction = "vse16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000???  :  Instruction = "vse32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000???  :  Instruction = "vse64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000???  :  Instruction = "vse8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000???  :  Instruction = "vse16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000???  :  Instruction = "vse32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000???  :  Instruction = "vse64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000???  :  Instruction = "vse8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000???  :  Instruction = "vse16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000???  :  Instruction = "vse32[ff].v,e16,mf2";
	    34'b0100111???????111?00111100?0000???  :  Instruction = "vse64[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000???  :  Instruction = "vse8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000???  :  Instruction = "vse16[ff].v,e16,m1";
	    34'b0100111???????110?00100000?0000???  :  Instruction = "vse32[ff].v,e16,m1";
	    34'b0100111???????111?00100000?0000???  :  Instruction = "vse64[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000???  :  Instruction = "vse8[ff].v,e16,m2";
	    34'b0100111???????101?00100100?0000???  :  Instruction = "vse16[ff].v,e16,m2";
	    34'b0100111???????110?00100100?0000???  :  Instruction = "vse32[ff].v,e16,m2";
	    34'b0100111???????111?00100100?0000???  :  Instruction = "vse64[ff].v,e16,m2";
	    34'b0100111???????000?00101000?0000???  :  Instruction = "vse8[ff].v,e16,m4";
	    34'b0100111???????101?00101000?0000???  :  Instruction = "vse16[ff].v,e16,m4";
	    34'b0100111???????110?00101000?0000???  :  Instruction = "vse32[ff].v,e16,m4";
	    34'b0100111???????000?00101100?0000???  :  Instruction = "vse8[ff].v,e16,m8";
	    34'b0100111???????101?00101100?0000???  :  Instruction = "vse16[ff].v,e16,m8";
	    34'b0100111???????000?001???0001000000  :  Instruction = "vs1r.v,e16";
	    34'b0100111???????101?00110110????????  :  Instruction = "vsse16.v,e16,mf8";
	    34'b0100111???????110?00110110????????  :  Instruction = "vsse32.v,e16,mf8";
	    34'b0100111???????111?00110110????????  :  Instruction = "vsse64.v,e16,mf8";
	    34'b0100111???????000?00111010????????  :  Instruction = "vsse8.v,e16,mf4";
	    34'b0100111???????101?00111010????????  :  Instruction = "vsse16.v,e16,mf4";
	    34'b0100111???????110?00111010????????  :  Instruction = "vsse32.v,e16,mf4";
	    34'b0100111???????111?00111010????????  :  Instruction = "vsse64.v,e16,mf4";
	    34'b0100111???????000?00111110????????  :  Instruction = "vsse8.v,e16,mf2";
	    34'b0100111???????101?00111110????????  :  Instruction = "vsse16.v,e16,mf2";
	    34'b0100111???????110?00111110????????  :  Instruction = "vsse32.v,e16,mf2";
	    34'b0100111???????111?00111110????????  :  Instruction = "vsse64.v,e16,mf2";
	    34'b0100111???????000?00100010????????  :  Instruction = "vsse8.v,e16,m1";
	    34'b0100111???????101?00100010????????  :  Instruction = "vsse16.v,e16,m1";
	    34'b0100111???????110?00100010????????  :  Instruction = "vsse32.v,e16,m1";
	    34'b0100111???????111?00100010????????  :  Instruction = "vsse64.v,e16,m1";
	    34'b0100111???????000?00100110????????  :  Instruction = "vsse8.v,e16,m2";
	    34'b0100111???????101?00100110????????  :  Instruction = "vsse16.v,e16,m2";
	    34'b0100111???????110?00100110????????  :  Instruction = "vsse32.v,e16,m2";
	    34'b0100111???????111?00100110????????  :  Instruction = "vsse64.v,e16,m2";
	    34'b0100111???????000?00101010????????  :  Instruction = "vsse8.v,e16,m4";
	    34'b0100111???????101?00101010????????  :  Instruction = "vsse16.v,e16,m4";
	    34'b0100111???????110?00101010????????  :  Instruction = "vsse32.v,e16,m4";
	    34'b0100111???????000?00101110????????  :  Instruction = "vsse8.v,e16,m8";
	    34'b0100111???????101?00101110????????  :  Instruction = "vsse16.v,e16,m8";
	    34'b0100111???????101?001101?1????????  :  Instruction = "vs[uo]xei16.v,e16,mf8";
	    34'b0100111???????110?001101?1????????  :  Instruction = "vs[uo]xei32.v,e16,mf8";
	    34'b0100111???????111?001101?1????????  :  Instruction = "vs[uo]xei64.v,e16,mf8";
	    34'b0100111???????000?001110?1????????  :  Instruction = "vs[uo]xei8.v,e16,mf4";
	    34'b0100111???????101?001110?1????????  :  Instruction = "vs[uo]xei16.v,e16,mf4";
	    34'b0100111???????110?001110?1????????  :  Instruction = "vs[uo]xei32.v,e16,mf4";
	    34'b0100111???????111?001110?1????????  :  Instruction = "vs[uo]xei64.v,e16,mf4";
	    34'b0100111???????000?001111?1????????  :  Instruction = "vs[uo]xei8.v,e16,mf2";
	    34'b0100111???????101?001111?1????????  :  Instruction = "vs[uo]xei16.v,e16,mf2";
	    34'b0100111???????110?001111?1????????  :  Instruction = "vs[uo]xei32.v,e16,mf2";
	    34'b0100111???????111?001111?1????????  :  Instruction = "vs[uo]xei64.v,e16,mf2";
	    34'b0100111???????000?001000?1????????  :  Instruction = "vs[uo]xei8.v,e16,m1";
	    34'b0100111???????101?001000?1????????  :  Instruction = "vs[uo]xei16.v,e16,m1";
	    34'b0100111???????110?001000?1????????  :  Instruction = "vs[uo]xei32.v,e16,m1";
	    34'b0100111???????111?001000?1????????  :  Instruction = "vs[uo]xei64.v,e16,m1";
	    34'b0100111???????000?001001?1????????  :  Instruction = "vs[uo]xei8.v,e16,m2";
	    34'b0100111???????101?001001?1????????  :  Instruction = "vs[uo]xei16.v,e16,m2";
	    34'b0100111???????110?001001?1????????  :  Instruction = "vs[uo]xei32.v,e16,m2";
	    34'b0100111???????111?001001?1????????  :  Instruction = "vs[uo]xei64.v,e16,m2";
	    34'b0100111???????000?001010?1????????  :  Instruction = "vs[uo]xei8.v,e16,m4";
	    34'b0100111???????101?001010?1????????  :  Instruction = "vs[uo]xei16.v,e16,m4";
	    34'b0100111???????110?001010?1????????  :  Instruction = "vs[uo]xei32.v,e16,m4";
	    34'b0100111???????000?001011?1????????  :  Instruction = "vs[uo]xei8.v,e16,m8";
	    34'b0100111???????101?001011?1????????  :  Instruction = "vs[uo]xei16.v,e16,m8";
	    34'b0100111???????101?00110100?0000001  :  Instruction = "vsseg2e16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000001  :  Instruction = "vsseg2e32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000001  :  Instruction = "vsseg2e64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000001  :  Instruction = "vsseg2e8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000001  :  Instruction = "vsseg2e16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000001  :  Instruction = "vsseg2e32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000001  :  Instruction = "vsseg2e64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000001  :  Instruction = "vsseg2e8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000001  :  Instruction = "vsseg2e16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000001  :  Instruction = "vsseg2e32[ff].v,e16,mf2";
	    34'b0100111???????111?00111100?0000001  :  Instruction = "vsseg2e64[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000001  :  Instruction = "vsseg2e8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000001  :  Instruction = "vsseg2e16[ff].v,e16,m1";
	    34'b0100111???????110?00100000?0000001  :  Instruction = "vsseg2e32[ff].v,e16,m1";
	    34'b0100111???????111?00100000?0000001  :  Instruction = "vsseg2e64[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000001  :  Instruction = "vsseg2e8[ff].v,e16,m2";
	    34'b0100111???????101?00100100?0000001  :  Instruction = "vsseg2e16[ff].v,e16,m2";
	    34'b0100111???????110?00100100?0000001  :  Instruction = "vsseg2e32[ff].v,e16,m2";
	    34'b0100111???????000?00101000?0000001  :  Instruction = "vsseg2e8[ff].v,e16,m4";
	    34'b0100111???????101?00101000?0000001  :  Instruction = "vsseg2e16[ff].v,e16,m4";
	    34'b0100111???????000?00101100?0000001  :  Instruction = "vsseg2e8[ff].v,e16,m8";
	    34'b0100111???????000?001???0001000001  :  Instruction = "vs2r.v,e16";
	    34'b0100111???????101?00110110?????001  :  Instruction = "vssseg2e16.v,e16,mf8";
	    34'b0100111???????110?00110110?????001  :  Instruction = "vssseg2e32.v,e16,mf8";
	    34'b0100111???????111?00110110?????001  :  Instruction = "vssseg2e64.v,e16,mf8";
	    34'b0100111???????000?00111010?????001  :  Instruction = "vssseg2e8.v,e16,mf4";
	    34'b0100111???????101?00111010?????001  :  Instruction = "vssseg2e16.v,e16,mf4";
	    34'b0100111???????110?00111010?????001  :  Instruction = "vssseg2e32.v,e16,mf4";
	    34'b0100111???????111?00111010?????001  :  Instruction = "vssseg2e64.v,e16,mf4";
	    34'b0100111???????000?00111110?????001  :  Instruction = "vssseg2e8.v,e16,mf2";
	    34'b0100111???????101?00111110?????001  :  Instruction = "vssseg2e16.v,e16,mf2";
	    34'b0100111???????110?00111110?????001  :  Instruction = "vssseg2e32.v,e16,mf2";
	    34'b0100111???????111?00111110?????001  :  Instruction = "vssseg2e64.v,e16,mf2";
	    34'b0100111???????000?00100010?????001  :  Instruction = "vssseg2e8.v,e16,m1";
	    34'b0100111???????101?00100010?????001  :  Instruction = "vssseg2e16.v,e16,m1";
	    34'b0100111???????110?00100010?????001  :  Instruction = "vssseg2e32.v,e16,m1";
	    34'b0100111???????111?00100010?????001  :  Instruction = "vssseg2e64.v,e16,m1";
	    34'b0100111???????000?00100110?????001  :  Instruction = "vssseg2e8.v,e16,m2";
	    34'b0100111???????101?00100110?????001  :  Instruction = "vssseg2e16.v,e16,m2";
	    34'b0100111???????110?00100110?????001  :  Instruction = "vssseg2e32.v,e16,m2";
	    34'b0100111???????000?00101010?????001  :  Instruction = "vssseg2e8.v,e16,m4";
	    34'b0100111???????101?00101010?????001  :  Instruction = "vssseg2e16.v,e16,m4";
	    34'b0100111???????000?00101110?????001  :  Instruction = "vssseg2e8.v,e16,m8";
	    34'b0100111???????101?001101?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e16,mf8";
	    34'b0100111???????110?001101?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e16,mf8";
	    34'b0100111???????111?001101?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e16,mf8";
	    34'b0100111???????000?001110?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e16,mf4";
	    34'b0100111???????101?001110?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e16,mf4";
	    34'b0100111???????110?001110?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e16,mf4";
	    34'b0100111???????111?001110?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e16,mf4";
	    34'b0100111???????000?001111?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e16,mf2";
	    34'b0100111???????101?001111?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e16,mf2";
	    34'b0100111???????110?001111?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e16,mf2";
	    34'b0100111???????111?001111?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e16,mf2";
	    34'b0100111???????000?001000?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e16,m1";
	    34'b0100111???????101?001000?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e16,m1";
	    34'b0100111???????110?001000?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e16,m1";
	    34'b0100111???????111?001000?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e16,m1";
	    34'b0100111???????000?001001?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e16,m2";
	    34'b0100111???????101?001001?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e16,m2";
	    34'b0100111???????110?001001?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e16,m2";
	    34'b0100111???????111?001001?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e16,m2";
	    34'b0100111???????000?001010?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e16,m4";
	    34'b0100111???????101?001010?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e16,m4";
	    34'b0100111???????110?001010?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e16,m4";
	    34'b0100111???????101?00110100?0000010  :  Instruction = "vsseg3e16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000010  :  Instruction = "vsseg3e32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000010  :  Instruction = "vsseg3e64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000010  :  Instruction = "vsseg3e8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000010  :  Instruction = "vsseg3e16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000010  :  Instruction = "vsseg3e32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000010  :  Instruction = "vsseg3e64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000010  :  Instruction = "vsseg3e8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000010  :  Instruction = "vsseg3e16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000010  :  Instruction = "vsseg3e32[ff].v,e16,mf2";
	    34'b0100111???????111?00111100?0000010  :  Instruction = "vsseg3e64[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000010  :  Instruction = "vsseg3e8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000010  :  Instruction = "vsseg3e16[ff].v,e16,m1";
	    34'b0100111???????110?00100000?0000010  :  Instruction = "vsseg3e32[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000010  :  Instruction = "vsseg3e8[ff].v,e16,m2";
	    34'b0100111???????101?00100100?0000010  :  Instruction = "vsseg3e16[ff].v,e16,m2";
	    34'b0100111???????000?00101000?0000010  :  Instruction = "vsseg3e8[ff].v,e16,m4";
	    34'b0100111???????101?00110110?????010  :  Instruction = "vssseg3e16.v,e16,mf8";
	    34'b0100111???????110?00110110?????010  :  Instruction = "vssseg3e32.v,e16,mf8";
	    34'b0100111???????111?00110110?????010  :  Instruction = "vssseg3e64.v,e16,mf8";
	    34'b0100111???????000?00111010?????010  :  Instruction = "vssseg3e8.v,e16,mf4";
	    34'b0100111???????101?00111010?????010  :  Instruction = "vssseg3e16.v,e16,mf4";
	    34'b0100111???????110?00111010?????010  :  Instruction = "vssseg3e32.v,e16,mf4";
	    34'b0100111???????111?00111010?????010  :  Instruction = "vssseg3e64.v,e16,mf4";
	    34'b0100111???????000?00111110?????010  :  Instruction = "vssseg3e8.v,e16,mf2";
	    34'b0100111???????101?00111110?????010  :  Instruction = "vssseg3e16.v,e16,mf2";
	    34'b0100111???????110?00111110?????010  :  Instruction = "vssseg3e32.v,e16,mf2";
	    34'b0100111???????111?00111110?????010  :  Instruction = "vssseg3e64.v,e16,mf2";
	    34'b0100111???????000?00100010?????010  :  Instruction = "vssseg3e8.v,e16,m1";
	    34'b0100111???????101?00100010?????010  :  Instruction = "vssseg3e16.v,e16,m1";
	    34'b0100111???????110?00100010?????010  :  Instruction = "vssseg3e32.v,e16,m1";
	    34'b0100111???????000?00100110?????010  :  Instruction = "vssseg3e8.v,e16,m2";
	    34'b0100111???????101?00100110?????010  :  Instruction = "vssseg3e16.v,e16,m2";
	    34'b0100111???????000?00101010?????010  :  Instruction = "vssseg3e8.v,e16,m4";
	    34'b0100111???????101?001101?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e16,mf8";
	    34'b0100111???????110?001101?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e16,mf8";
	    34'b0100111???????111?001101?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e16,mf8";
	    34'b0100111???????000?001110?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e16,mf4";
	    34'b0100111???????101?001110?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e16,mf4";
	    34'b0100111???????110?001110?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e16,mf4";
	    34'b0100111???????111?001110?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e16,mf4";
	    34'b0100111???????000?001111?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e16,mf2";
	    34'b0100111???????101?001111?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e16,mf2";
	    34'b0100111???????110?001111?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e16,mf2";
	    34'b0100111???????111?001111?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e16,mf2";
	    34'b0100111???????000?001000?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e16,m1";
	    34'b0100111???????101?001000?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e16,m1";
	    34'b0100111???????110?001000?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e16,m1";
	    34'b0100111???????111?001000?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e16,m1";
	    34'b0100111???????000?001001?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e16,m2";
	    34'b0100111???????101?001001?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e16,m2";
	    34'b0100111???????110?001001?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e16,m2";
	    34'b0100111???????111?001001?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e16,m2";
	    34'b0100111???????101?00110100?0000011  :  Instruction = "vsseg4e16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000011  :  Instruction = "vsseg4e32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000011  :  Instruction = "vsseg4e64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000011  :  Instruction = "vsseg4e8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000011  :  Instruction = "vsseg4e16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000011  :  Instruction = "vsseg4e32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000011  :  Instruction = "vsseg4e64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000011  :  Instruction = "vsseg4e8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000011  :  Instruction = "vsseg4e16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000011  :  Instruction = "vsseg4e32[ff].v,e16,mf2";
	    34'b0100111???????111?00111100?0000011  :  Instruction = "vsseg4e64[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000011  :  Instruction = "vsseg4e8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000011  :  Instruction = "vsseg4e16[ff].v,e16,m1";
	    34'b0100111???????110?00100000?0000011  :  Instruction = "vsseg4e32[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000011  :  Instruction = "vsseg4e8[ff].v,e16,m2";
	    34'b0100111???????101?00100100?0000011  :  Instruction = "vsseg4e16[ff].v,e16,m2";
	    34'b0100111???????000?00101000?0000011  :  Instruction = "vsseg4e8[ff].v,e16,m4";
	    34'b0100111???????101?00110110?????011  :  Instruction = "vssseg4e16.v,e16,mf8";
	    34'b0100111???????110?00110110?????011  :  Instruction = "vssseg4e32.v,e16,mf8";
	    34'b0100111???????111?00110110?????011  :  Instruction = "vssseg4e64.v,e16,mf8";
	    34'b0100111???????000?00111010?????011  :  Instruction = "vssseg4e8.v,e16,mf4";
	    34'b0100111???????101?00111010?????011  :  Instruction = "vssseg4e16.v,e16,mf4";
	    34'b0100111???????110?00111010?????011  :  Instruction = "vssseg4e32.v,e16,mf4";
	    34'b0100111???????111?00111010?????011  :  Instruction = "vssseg4e64.v,e16,mf4";
	    34'b0100111???????000?00111110?????011  :  Instruction = "vssseg4e8.v,e16,mf2";
	    34'b0100111???????101?00111110?????011  :  Instruction = "vssseg4e16.v,e16,mf2";
	    34'b0100111???????110?00111110?????011  :  Instruction = "vssseg4e32.v,e16,mf2";
	    34'b0100111???????111?00111110?????011  :  Instruction = "vssseg4e64.v,e16,mf2";
	    34'b0100111???????000?00100010?????011  :  Instruction = "vssseg4e8.v,e16,m1";
	    34'b0100111???????101?00100010?????011  :  Instruction = "vssseg4e16.v,e16,m1";
	    34'b0100111???????110?00100010?????011  :  Instruction = "vssseg4e32.v,e16,m1";
	    34'b0100111???????000?00100110?????011  :  Instruction = "vssseg4e8.v,e16,m2";
	    34'b0100111???????101?00100110?????011  :  Instruction = "vssseg4e16.v,e16,m2";
	    34'b0100111???????000?00101010?????011  :  Instruction = "vssseg4e8.v,e16,m4";
	    34'b0100111???????000?001???0001000011  :  Instruction = "vs4r.v,e16";
	    34'b0100111???????101?001101?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e16,mf8";
	    34'b0100111???????110?001101?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e16,mf8";
	    34'b0100111???????111?001101?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e16,mf8";
	    34'b0100111???????000?001110?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e16,mf4";
	    34'b0100111???????101?001110?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e16,mf4";
	    34'b0100111???????110?001110?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e16,mf4";
	    34'b0100111???????111?001110?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e16,mf4";
	    34'b0100111???????000?001111?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e16,mf2";
	    34'b0100111???????101?001111?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e16,mf2";
	    34'b0100111???????110?001111?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e16,mf2";
	    34'b0100111???????111?001111?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e16,mf2";
	    34'b0100111???????000?001000?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e16,m1";
	    34'b0100111???????101?001000?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e16,m1";
	    34'b0100111???????110?001000?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e16,m1";
	    34'b0100111???????111?001000?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e16,m1";
	    34'b0100111???????000?001001?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e16,m2";
	    34'b0100111???????101?001001?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e16,m2";
	    34'b0100111???????110?001001?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e16,m2";
	    34'b0100111???????111?001001?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e16,m2";
	    34'b0100111???????101?00110100?0000100  :  Instruction = "vsseg5e16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000100  :  Instruction = "vsseg5e32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000100  :  Instruction = "vsseg5e64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000100  :  Instruction = "vsseg5e8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000100  :  Instruction = "vsseg5e16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000100  :  Instruction = "vsseg5e32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000100  :  Instruction = "vsseg5e64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000100  :  Instruction = "vsseg5e8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000100  :  Instruction = "vsseg5e16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000100  :  Instruction = "vsseg5e32[ff].v,e16,mf2";
	    34'b0100111???????111?00111100?0000100  :  Instruction = "vsseg5e64[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000100  :  Instruction = "vsseg5e8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000100  :  Instruction = "vsseg5e16[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000100  :  Instruction = "vsseg5e8[ff].v,e16,m2";
	    34'b0100111???????101?00110110?????100  :  Instruction = "vssseg5e16.v,e16,mf8";
	    34'b0100111???????110?00110110?????100  :  Instruction = "vssseg5e32.v,e16,mf8";
	    34'b0100111???????111?00110110?????100  :  Instruction = "vssseg5e64.v,e16,mf8";
	    34'b0100111???????000?00111010?????100  :  Instruction = "vssseg5e8.v,e16,mf4";
	    34'b0100111???????101?00111010?????100  :  Instruction = "vssseg5e16.v,e16,mf4";
	    34'b0100111???????110?00111010?????100  :  Instruction = "vssseg5e32.v,e16,mf4";
	    34'b0100111???????111?00111010?????100  :  Instruction = "vssseg5e64.v,e16,mf4";
	    34'b0100111???????000?00111110?????100  :  Instruction = "vssseg5e8.v,e16,mf2";
	    34'b0100111???????101?00111110?????100  :  Instruction = "vssseg5e16.v,e16,mf2";
	    34'b0100111???????110?00111110?????100  :  Instruction = "vssseg5e32.v,e16,mf2";
	    34'b0100111???????000?00100010?????100  :  Instruction = "vssseg5e8.v,e16,m1";
	    34'b0100111???????101?00100010?????100  :  Instruction = "vssseg5e16.v,e16,m1";
	    34'b0100111???????000?00100110?????100  :  Instruction = "vssseg5e8.v,e16,m2";
	    34'b0100111???????101?001101?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e16,mf8";
	    34'b0100111???????110?001101?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e16,mf8";
	    34'b0100111???????111?001101?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e16,mf8";
	    34'b0100111???????000?001110?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e16,mf4";
	    34'b0100111???????101?001110?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e16,mf4";
	    34'b0100111???????110?001110?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e16,mf4";
	    34'b0100111???????111?001110?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e16,mf4";
	    34'b0100111???????000?001111?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e16,mf2";
	    34'b0100111???????101?001111?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e16,mf2";
	    34'b0100111???????110?001111?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e16,mf2";
	    34'b0100111???????111?001111?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e16,mf2";
	    34'b0100111???????000?001000?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e16,m1";
	    34'b0100111???????101?001000?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e16,m1";
	    34'b0100111???????110?001000?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e16,m1";
	    34'b0100111???????111?001000?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e16,m1";
	    34'b0100111???????101?00110100?0000101  :  Instruction = "vsseg6e16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000101  :  Instruction = "vsseg6e32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000101  :  Instruction = "vsseg6e64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000101  :  Instruction = "vsseg6e8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000101  :  Instruction = "vsseg6e16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000101  :  Instruction = "vsseg6e32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000101  :  Instruction = "vsseg6e64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000101  :  Instruction = "vsseg6e8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000101  :  Instruction = "vsseg6e16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000101  :  Instruction = "vsseg6e32[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000101  :  Instruction = "vsseg6e8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000101  :  Instruction = "vsseg6e16[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000101  :  Instruction = "vsseg6e8[ff].v,e16,m2";
	    34'b0100111???????101?00110110?????101  :  Instruction = "vssseg6e16.v,e16,mf8";
	    34'b0100111???????110?00110110?????101  :  Instruction = "vssseg6e32.v,e16,mf8";
	    34'b0100111???????111?00110110?????101  :  Instruction = "vssseg6e64.v,e16,mf8";
	    34'b0100111???????000?00111010?????101  :  Instruction = "vssseg6e8.v,e16,mf4";
	    34'b0100111???????101?00111010?????101  :  Instruction = "vssseg6e16.v,e16,mf4";
	    34'b0100111???????110?00111010?????101  :  Instruction = "vssseg6e32.v,e16,mf4";
	    34'b0100111???????111?00111010?????101  :  Instruction = "vssseg6e64.v,e16,mf4";
	    34'b0100111???????000?00111110?????101  :  Instruction = "vssseg6e8.v,e16,mf2";
	    34'b0100111???????101?00111110?????101  :  Instruction = "vssseg6e16.v,e16,mf2";
	    34'b0100111???????110?00111110?????101  :  Instruction = "vssseg6e32.v,e16,mf2";
	    34'b0100111???????000?00100010?????101  :  Instruction = "vssseg6e8.v,e16,m1";
	    34'b0100111???????101?00100010?????101  :  Instruction = "vssseg6e16.v,e16,m1";
	    34'b0100111???????000?00100110?????101  :  Instruction = "vssseg6e8.v,e16,m2";
	    34'b0100111???????101?001101?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e16,mf8";
	    34'b0100111???????110?001101?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e16,mf8";
	    34'b0100111???????111?001101?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e16,mf8";
	    34'b0100111???????000?001110?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e16,mf4";
	    34'b0100111???????101?001110?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e16,mf4";
	    34'b0100111???????110?001110?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e16,mf4";
	    34'b0100111???????111?001110?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e16,mf4";
	    34'b0100111???????000?001111?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e16,mf2";
	    34'b0100111???????101?001111?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e16,mf2";
	    34'b0100111???????110?001111?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e16,mf2";
	    34'b0100111???????111?001111?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e16,mf2";
	    34'b0100111???????000?001000?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e16,m1";
	    34'b0100111???????101?001000?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e16,m1";
	    34'b0100111???????110?001000?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e16,m1";
	    34'b0100111???????111?001000?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e16,m1";
	    34'b0100111???????101?00110100?0000110  :  Instruction = "vsseg7e16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000110  :  Instruction = "vsseg7e32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000110  :  Instruction = "vsseg7e64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000110  :  Instruction = "vsseg7e8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000110  :  Instruction = "vsseg7e16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000110  :  Instruction = "vsseg7e32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000110  :  Instruction = "vsseg7e64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000110  :  Instruction = "vsseg7e8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000110  :  Instruction = "vsseg7e16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000110  :  Instruction = "vsseg7e32[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000110  :  Instruction = "vsseg7e8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000110  :  Instruction = "vsseg7e16[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000110  :  Instruction = "vsseg7e8[ff].v,e16,m2";
	    34'b0100111???????101?00110110?????110  :  Instruction = "vssseg7e16.v,e16,mf8";
	    34'b0100111???????110?00110110?????110  :  Instruction = "vssseg7e32.v,e16,mf8";
	    34'b0100111???????111?00110110?????110  :  Instruction = "vssseg7e64.v,e16,mf8";
	    34'b0100111???????000?00111010?????110  :  Instruction = "vssseg7e8.v,e16,mf4";
	    34'b0100111???????101?00111010?????110  :  Instruction = "vssseg7e16.v,e16,mf4";
	    34'b0100111???????110?00111010?????110  :  Instruction = "vssseg7e32.v,e16,mf4";
	    34'b0100111???????111?00111010?????110  :  Instruction = "vssseg7e64.v,e16,mf4";
	    34'b0100111???????000?00111110?????110  :  Instruction = "vssseg7e8.v,e16,mf2";
	    34'b0100111???????101?00111110?????110  :  Instruction = "vssseg7e16.v,e16,mf2";
	    34'b0100111???????110?00111110?????110  :  Instruction = "vssseg7e32.v,e16,mf2";
	    34'b0100111???????000?00100010?????110  :  Instruction = "vssseg7e8.v,e16,m1";
	    34'b0100111???????101?00100010?????110  :  Instruction = "vssseg7e16.v,e16,m1";
	    34'b0100111???????000?00100110?????110  :  Instruction = "vssseg7e8.v,e16,m2";
	    34'b0100111???????101?001101?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e16,mf8";
	    34'b0100111???????110?001101?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e16,mf8";
	    34'b0100111???????111?001101?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e16,mf8";
	    34'b0100111???????000?001110?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e16,mf4";
	    34'b0100111???????101?001110?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e16,mf4";
	    34'b0100111???????110?001110?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e16,mf4";
	    34'b0100111???????111?001110?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e16,mf4";
	    34'b0100111???????000?001111?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e16,mf2";
	    34'b0100111???????101?001111?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e16,mf2";
	    34'b0100111???????110?001111?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e16,mf2";
	    34'b0100111???????111?001111?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e16,mf2";
	    34'b0100111???????000?001000?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e16,m1";
	    34'b0100111???????101?001000?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e16,m1";
	    34'b0100111???????110?001000?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e16,m1";
	    34'b0100111???????111?001000?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e16,m1";
	    34'b0100111???????101?00110100?0000111  :  Instruction = "vsseg8e16[ff].v,e16,mf8";
	    34'b0100111???????110?00110100?0000111  :  Instruction = "vsseg8e32[ff].v,e16,mf8";
	    34'b0100111???????111?00110100?0000111  :  Instruction = "vsseg8e64[ff].v,e16,mf8";
	    34'b0100111???????000?00111000?0000111  :  Instruction = "vsseg8e8[ff].v,e16,mf4";
	    34'b0100111???????101?00111000?0000111  :  Instruction = "vsseg8e16[ff].v,e16,mf4";
	    34'b0100111???????110?00111000?0000111  :  Instruction = "vsseg8e32[ff].v,e16,mf4";
	    34'b0100111???????111?00111000?0000111  :  Instruction = "vsseg8e64[ff].v,e16,mf4";
	    34'b0100111???????000?00111100?0000111  :  Instruction = "vsseg8e8[ff].v,e16,mf2";
	    34'b0100111???????101?00111100?0000111  :  Instruction = "vsseg8e16[ff].v,e16,mf2";
	    34'b0100111???????110?00111100?0000111  :  Instruction = "vsseg8e32[ff].v,e16,mf2";
	    34'b0100111???????000?00100000?0000111  :  Instruction = "vsseg8e8[ff].v,e16,m1";
	    34'b0100111???????101?00100000?0000111  :  Instruction = "vsseg8e16[ff].v,e16,m1";
	    34'b0100111???????000?00100100?0000111  :  Instruction = "vsseg8e8[ff].v,e16,m2";
	    34'b0100111???????000?001???0001000111  :  Instruction = "vs8r.v,e16";
	    34'b0100111???????101?00110110?????111  :  Instruction = "vssseg8e16.v,e16,mf8";
	    34'b0100111???????110?00110110?????111  :  Instruction = "vssseg8e32.v,e16,mf8";
	    34'b0100111???????111?00110110?????111  :  Instruction = "vssseg8e64.v,e16,mf8";
	    34'b0100111???????000?00111010?????111  :  Instruction = "vssseg8e8.v,e16,mf4";
	    34'b0100111???????101?00111010?????111  :  Instruction = "vssseg8e16.v,e16,mf4";
	    34'b0100111???????110?00111010?????111  :  Instruction = "vssseg8e32.v,e16,mf4";
	    34'b0100111???????111?00111010?????111  :  Instruction = "vssseg8e64.v,e16,mf4";
	    34'b0100111???????000?00111110?????111  :  Instruction = "vssseg8e8.v,e16,mf2";
	    34'b0100111???????101?00111110?????111  :  Instruction = "vssseg8e16.v,e16,mf2";
	    34'b0100111???????110?00111110?????111  :  Instruction = "vssseg8e32.v,e16,mf2";
	    34'b0100111???????000?00100010?????111  :  Instruction = "vssseg8e8.v,e16,m1";
	    34'b0100111???????101?00100010?????111  :  Instruction = "vssseg8e16.v,e16,m1";
	    34'b0100111???????000?00100110?????111  :  Instruction = "vssseg8e8.v,e16,m2";
	    34'b0100111???????101?001101?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e16,mf8";
	    34'b0100111???????110?001101?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e16,mf8";
	    34'b0100111???????111?001101?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e16,mf8";
	    34'b0100111???????000?001110?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e16,mf4";
	    34'b0100111???????101?001110?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e16,mf4";
	    34'b0100111???????110?001110?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e16,mf4";
	    34'b0100111???????111?001110?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e16,mf4";
	    34'b0100111???????000?001111?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e16,mf2";
	    34'b0100111???????101?001111?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e16,mf2";
	    34'b0100111???????110?001111?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e16,mf2";
	    34'b0100111???????111?001111?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e16,mf2";
	    34'b0100111???????000?001000?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e16,m1";
	    34'b0100111???????101?001000?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e16,m1";
	    34'b0100111???????110?001000?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e16,m1";
	    34'b0100111???????111?001000?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e16,m1";
	    34'b0000111???????110?01010100?0000???  :  Instruction = "vle32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000???  :  Instruction = "vle64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000???  :  Instruction = "vle16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000???  :  Instruction = "vle32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000???  :  Instruction = "vle64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000???  :  Instruction = "vle8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000???  :  Instruction = "vle16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000???  :  Instruction = "vle32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000???  :  Instruction = "vle64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000???  :  Instruction = "vle8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000???  :  Instruction = "vle16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000???  :  Instruction = "vle32[ff].v,e32,m1";
	    34'b0000111???????111?01000000?0000???  :  Instruction = "vle64[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000???  :  Instruction = "vle8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000???  :  Instruction = "vle16[ff].v,e32,m2";
	    34'b0000111???????110?01000100?0000???  :  Instruction = "vle32[ff].v,e32,m2";
	    34'b0000111???????111?01000100?0000???  :  Instruction = "vle64[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000???  :  Instruction = "vle8[ff].v,e32,m4";
	    34'b0000111???????101?01001000?0000???  :  Instruction = "vle16[ff].v,e32,m4";
	    34'b0000111???????110?01001000?0000???  :  Instruction = "vle32[ff].v,e32,m4";
	    34'b0000111???????111?01001000?0000???  :  Instruction = "vle64[ff].v,e32,m4";
	    34'b0000111???????000?01001100?0000???  :  Instruction = "vle8[ff].v,e32,m8";
	    34'b0000111???????101?01001100?0000???  :  Instruction = "vle16[ff].v,e32,m8";
	    34'b0000111???????110?01001100?0000???  :  Instruction = "vle32[ff].v,e32,m8";
	    34'b0000111???????000?010???0001000000  :  Instruction = "vl1re8.v,e32";
	    34'b0000111???????101?010???0001000000  :  Instruction = "vl1re16.v,e32";
	    34'b0000111???????110?010???0001000000  :  Instruction = "vl1re32.v,e32";
	    34'b0000111???????111?010???0001000000  :  Instruction = "vl1re64.v,e32";
	    34'b0000111???????110?01010110????????  :  Instruction = "vlse32.v,e32,mf8";
	    34'b0000111???????111?01010110????????  :  Instruction = "vlse64.v,e32,mf8";
	    34'b0000111???????101?01011010????????  :  Instruction = "vlse16.v,e32,mf4";
	    34'b0000111???????110?01011010????????  :  Instruction = "vlse32.v,e32,mf4";
	    34'b0000111???????111?01011010????????  :  Instruction = "vlse64.v,e32,mf4";
	    34'b0000111???????000?01011110????????  :  Instruction = "vlse8.v,e32,mf2";
	    34'b0000111???????101?01011110????????  :  Instruction = "vlse16.v,e32,mf2";
	    34'b0000111???????110?01011110????????  :  Instruction = "vlse32.v,e32,mf2";
	    34'b0000111???????111?01011110????????  :  Instruction = "vlse64.v,e32,mf2";
	    34'b0000111???????000?01000010????????  :  Instruction = "vlse8.v,e32,m1";
	    34'b0000111???????101?01000010????????  :  Instruction = "vlse16.v,e32,m1";
	    34'b0000111???????110?01000010????????  :  Instruction = "vlse32.v,e32,m1";
	    34'b0000111???????111?01000010????????  :  Instruction = "vlse64.v,e32,m1";
	    34'b0000111???????000?01000110????????  :  Instruction = "vlse8.v,e32,m2";
	    34'b0000111???????101?01000110????????  :  Instruction = "vlse16.v,e32,m2";
	    34'b0000111???????110?01000110????????  :  Instruction = "vlse32.v,e32,m2";
	    34'b0000111???????111?01000110????????  :  Instruction = "vlse64.v,e32,m2";
	    34'b0000111???????000?01001010????????  :  Instruction = "vlse8.v,e32,m4";
	    34'b0000111???????101?01001010????????  :  Instruction = "vlse16.v,e32,m4";
	    34'b0000111???????110?01001010????????  :  Instruction = "vlse32.v,e32,m4";
	    34'b0000111???????111?01001010????????  :  Instruction = "vlse64.v,e32,m4";
	    34'b0000111???????000?01001110????????  :  Instruction = "vlse8.v,e32,m8";
	    34'b0000111???????101?01001110????????  :  Instruction = "vlse16.v,e32,m8";
	    34'b0000111???????110?01001110????????  :  Instruction = "vlse32.v,e32,m8";
	    34'b0000111???????110?010101?1????????  :  Instruction = "vl[uo]xei32.v,e32,mf8";
	    34'b0000111???????111?010101?1????????  :  Instruction = "vl[uo]xei64.v,e32,mf8";
	    34'b0000111???????101?010110?1????????  :  Instruction = "vl[uo]xei16.v,e32,mf4";
	    34'b0000111???????110?010110?1????????  :  Instruction = "vl[uo]xei32.v,e32,mf4";
	    34'b0000111???????111?010110?1????????  :  Instruction = "vl[uo]xei64.v,e32,mf4";
	    34'b0000111???????000?010111?1????????  :  Instruction = "vl[uo]xei8.v,e32,mf2";
	    34'b0000111???????101?010111?1????????  :  Instruction = "vl[uo]xei16.v,e32,mf2";
	    34'b0000111???????110?010111?1????????  :  Instruction = "vl[uo]xei32.v,e32,mf2";
	    34'b0000111???????111?010111?1????????  :  Instruction = "vl[uo]xei64.v,e32,mf2";
	    34'b0000111???????000?010000?1????????  :  Instruction = "vl[uo]xei8.v,e32,m1";
	    34'b0000111???????101?010000?1????????  :  Instruction = "vl[uo]xei16.v,e32,m1";
	    34'b0000111???????110?010000?1????????  :  Instruction = "vl[uo]xei32.v,e32,m1";
	    34'b0000111???????111?010000?1????????  :  Instruction = "vl[uo]xei64.v,e32,m1";
	    34'b0000111???????000?010001?1????????  :  Instruction = "vl[uo]xei8.v,e32,m2";
	    34'b0000111???????101?010001?1????????  :  Instruction = "vl[uo]xei16.v,e32,m2";
	    34'b0000111???????110?010001?1????????  :  Instruction = "vl[uo]xei32.v,e32,m2";
	    34'b0000111???????111?010001?1????????  :  Instruction = "vl[uo]xei64.v,e32,m2";
	    34'b0000111???????000?010010?1????????  :  Instruction = "vl[uo]xei8.v,e32,m4";
	    34'b0000111???????101?010010?1????????  :  Instruction = "vl[uo]xei16.v,e32,m4";
	    34'b0000111???????110?010010?1????????  :  Instruction = "vl[uo]xei32.v,e32,m4";
	    34'b0000111???????111?010010?1????????  :  Instruction = "vl[uo]xei64.v,e32,m4";
	    34'b0000111???????000?010011?1????????  :  Instruction = "vl[uo]xei8.v,e32,m8";
	    34'b0000111???????101?010011?1????????  :  Instruction = "vl[uo]xei16.v,e32,m8";
	    34'b0000111???????110?010011?1????????  :  Instruction = "vl[uo]xei32.v,e32,m8";
	    34'b0000111???????110?01010100?0000001  :  Instruction = "vlseg2e32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000001  :  Instruction = "vlseg2e64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000001  :  Instruction = "vlseg2e16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000001  :  Instruction = "vlseg2e32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000001  :  Instruction = "vlseg2e64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000001  :  Instruction = "vlseg2e8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000001  :  Instruction = "vlseg2e16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000001  :  Instruction = "vlseg2e32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000001  :  Instruction = "vlseg2e64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000001  :  Instruction = "vlseg2e8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000001  :  Instruction = "vlseg2e16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000001  :  Instruction = "vlseg2e32[ff].v,e32,m1";
	    34'b0000111???????111?01000000?0000001  :  Instruction = "vlseg2e64[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000001  :  Instruction = "vlseg2e8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000001  :  Instruction = "vlseg2e16[ff].v,e32,m2";
	    34'b0000111???????110?01000100?0000001  :  Instruction = "vlseg2e32[ff].v,e32,m2";
	    34'b0000111???????111?01000100?0000001  :  Instruction = "vlseg2e64[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000001  :  Instruction = "vlseg2e8[ff].v,e32,m4";
	    34'b0000111???????101?01001000?0000001  :  Instruction = "vlseg2e16[ff].v,e32,m4";
	    34'b0000111???????110?01001000?0000001  :  Instruction = "vlseg2e32[ff].v,e32,m4";
	    34'b0000111???????000?01001100?0000001  :  Instruction = "vlseg2e8[ff].v,e32,m8";
	    34'b0000111???????101?01001100?0000001  :  Instruction = "vlseg2e16[ff].v,e32,m8";
	    34'b0000111???????111?01001100?0000001  :  Instruction = "vlseg2e64[ff].v,e32,m8";
	    34'b0000111???????000?010???0001000001  :  Instruction = "vl2re8.v,e32";
	    34'b0000111???????101?010???0001000001  :  Instruction = "vl2re16.v,e32";
	    34'b0000111???????110?010???0001000001  :  Instruction = "vl2re32.v,e32";
	    34'b0000111???????111?010???0001000001  :  Instruction = "vl2re64.v,e32";
	    34'b0000111???????110?01010110?????001  :  Instruction = "vlsseg2e32.v,e32,mf8";
	    34'b0000111???????111?01010110?????001  :  Instruction = "vlsseg2e64.v,e32,mf8";
	    34'b0000111???????101?01011010?????001  :  Instruction = "vlsseg2e16.v,e32,mf4";
	    34'b0000111???????110?01011010?????001  :  Instruction = "vlsseg2e32.v,e32,mf4";
	    34'b0000111???????111?01011010?????001  :  Instruction = "vlsseg2e64.v,e32,mf4";
	    34'b0000111???????000?01011110?????001  :  Instruction = "vlsseg2e8.v,e32,mf2";
	    34'b0000111???????101?01011110?????001  :  Instruction = "vlsseg2e16.v,e32,mf2";
	    34'b0000111???????110?01011110?????001  :  Instruction = "vlsseg2e32.v,e32,mf2";
	    34'b0000111???????111?01011110?????001  :  Instruction = "vlsseg2e64.v,e32,mf2";
	    34'b0000111???????000?01000010?????001  :  Instruction = "vlsseg2e8.v,e32,m1";
	    34'b0000111???????101?01000010?????001  :  Instruction = "vlsseg2e16.v,e32,m1";
	    34'b0000111???????110?01000010?????001  :  Instruction = "vlsseg2e32.v,e32,m1";
	    34'b0000111???????111?01000010?????001  :  Instruction = "vlsseg2e64.v,e32,m1";
	    34'b0000111???????000?01000110?????001  :  Instruction = "vlsseg2e8.v,e32,m2";
	    34'b0000111???????101?01000110?????001  :  Instruction = "vlsseg2e16.v,e32,m2";
	    34'b0000111???????110?01000110?????001  :  Instruction = "vlsseg2e32.v,e32,m2";
	    34'b0000111???????111?01000110?????001  :  Instruction = "vlsseg2e64.v,e32,m2";
	    34'b0000111???????000?01001010?????001  :  Instruction = "vlsseg2e8.v,e32,m4";
	    34'b0000111???????101?01001010?????001  :  Instruction = "vlsseg2e16.v,e32,m4";
	    34'b0000111???????110?01001010?????001  :  Instruction = "vlsseg2e32.v,e32,m4";
	    34'b0000111???????000?01001110?????001  :  Instruction = "vlsseg2e8.v,e32,m8";
	    34'b0000111???????101?01001110?????001  :  Instruction = "vlsseg2e16.v,e32,m8";
	    34'b0000111???????110?010101?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e32,mf8";
	    34'b0000111???????111?010101?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e32,mf8";
	    34'b0000111???????101?010110?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e32,mf4";
	    34'b0000111???????110?010110?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e32,mf4";
	    34'b0000111???????111?010110?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e32,mf4";
	    34'b0000111???????000?010111?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e32,mf2";
	    34'b0000111???????101?010111?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e32,mf2";
	    34'b0000111???????110?010111?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e32,mf2";
	    34'b0000111???????111?010111?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e32,mf2";
	    34'b0000111???????000?010000?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e32,m1";
	    34'b0000111???????101?010000?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e32,m1";
	    34'b0000111???????110?010000?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e32,m1";
	    34'b0000111???????111?010000?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e32,m1";
	    34'b0000111???????000?010001?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e32,m2";
	    34'b0000111???????101?010001?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e32,m2";
	    34'b0000111???????110?010001?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e32,m2";
	    34'b0000111???????111?010001?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e32,m2";
	    34'b0000111???????000?010010?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e32,m4";
	    34'b0000111???????101?010010?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e32,m4";
	    34'b0000111???????110?010010?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e32,m4";
	    34'b0000111???????111?010010?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e32,m4";
	    34'b0000111???????110?01010100?0000010  :  Instruction = "vlseg3e32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000010  :  Instruction = "vlseg3e64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000010  :  Instruction = "vlseg3e16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000010  :  Instruction = "vlseg3e32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000010  :  Instruction = "vlseg3e64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000010  :  Instruction = "vlseg3e8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000010  :  Instruction = "vlseg3e16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000010  :  Instruction = "vlseg3e32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000010  :  Instruction = "vlseg3e64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000010  :  Instruction = "vlseg3e8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000010  :  Instruction = "vlseg3e16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000010  :  Instruction = "vlseg3e32[ff].v,e32,m1";
	    34'b0000111???????111?01000000?0000010  :  Instruction = "vlseg3e64[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000010  :  Instruction = "vlseg3e8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000010  :  Instruction = "vlseg3e16[ff].v,e32,m2";
	    34'b0000111???????110?01000100?0000010  :  Instruction = "vlseg3e32[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000010  :  Instruction = "vlseg3e8[ff].v,e32,m4";
	    34'b0000111???????101?01001000?0000010  :  Instruction = "vlseg3e16[ff].v,e32,m4";
	    34'b0000111???????000?01001100?0000010  :  Instruction = "vlseg3e8[ff].v,e32,m8";
	    34'b0000111???????110?01010110?????010  :  Instruction = "vlsseg3e32.v,e32,mf8";
	    34'b0000111???????111?01010110?????010  :  Instruction = "vlsseg3e64.v,e32,mf8";
	    34'b0000111???????101?01011010?????010  :  Instruction = "vlsseg3e16.v,e32,mf4";
	    34'b0000111???????110?01011010?????010  :  Instruction = "vlsseg3e32.v,e32,mf4";
	    34'b0000111???????111?01011010?????010  :  Instruction = "vlsseg3e64.v,e32,mf4";
	    34'b0000111???????000?01011110?????010  :  Instruction = "vlsseg3e8.v,e32,mf2";
	    34'b0000111???????101?01011110?????010  :  Instruction = "vlsseg3e16.v,e32,mf2";
	    34'b0000111???????110?01011110?????010  :  Instruction = "vlsseg3e32.v,e32,mf2";
	    34'b0000111???????111?01011110?????010  :  Instruction = "vlsseg3e64.v,e32,mf2";
	    34'b0000111???????000?01000010?????010  :  Instruction = "vlsseg3e8.v,e32,m1";
	    34'b0000111???????101?01000010?????010  :  Instruction = "vlsseg3e16.v,e32,m1";
	    34'b0000111???????110?01000010?????010  :  Instruction = "vlsseg3e32.v,e32,m1";
	    34'b0000111???????111?01000010?????010  :  Instruction = "vlsseg3e64.v,e32,m1";
	    34'b0000111???????000?01000110?????010  :  Instruction = "vlsseg3e8.v,e32,m2";
	    34'b0000111???????101?01000110?????010  :  Instruction = "vlsseg3e16.v,e32,m2";
	    34'b0000111???????110?01000110?????010  :  Instruction = "vlsseg3e32.v,e32,m2";
	    34'b0000111???????000?01001010?????010  :  Instruction = "vlsseg3e8.v,e32,m4";
	    34'b0000111???????101?01001010?????010  :  Instruction = "vlsseg3e16.v,e32,m4";
	    34'b0000111???????000?01001110?????010  :  Instruction = "vlsseg3e8.v,e32,m8";
	    34'b0000111???????110?010101?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e32,mf8";
	    34'b0000111???????111?010101?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e32,mf8";
	    34'b0000111???????101?010110?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e32,mf4";
	    34'b0000111???????110?010110?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e32,mf4";
	    34'b0000111???????111?010110?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e32,mf4";
	    34'b0000111???????000?010111?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e32,mf2";
	    34'b0000111???????101?010111?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e32,mf2";
	    34'b0000111???????110?010111?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e32,mf2";
	    34'b0000111???????111?010111?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e32,mf2";
	    34'b0000111???????000?010000?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e32,m1";
	    34'b0000111???????101?010000?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e32,m1";
	    34'b0000111???????110?010000?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e32,m1";
	    34'b0000111???????111?010000?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e32,m1";
	    34'b0000111???????000?010001?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e32,m2";
	    34'b0000111???????101?010001?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e32,m2";
	    34'b0000111???????110?010001?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e32,m2";
	    34'b0000111???????111?010001?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e32,m2";
	    34'b0000111???????110?01010100?0000011  :  Instruction = "vlseg4e32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000011  :  Instruction = "vlseg4e64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000011  :  Instruction = "vlseg4e16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000011  :  Instruction = "vlseg4e32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000011  :  Instruction = "vlseg4e64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000011  :  Instruction = "vlseg4e8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000011  :  Instruction = "vlseg4e16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000011  :  Instruction = "vlseg4e32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000011  :  Instruction = "vlseg4e64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000011  :  Instruction = "vlseg4e8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000011  :  Instruction = "vlseg4e16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000011  :  Instruction = "vlseg4e32[ff].v,e32,m1";
	    34'b0000111???????111?01000000?0000011  :  Instruction = "vlseg4e64[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000011  :  Instruction = "vlseg4e8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000011  :  Instruction = "vlseg4e16[ff].v,e32,m2";
	    34'b0000111???????110?01000100?0000011  :  Instruction = "vlseg4e32[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000011  :  Instruction = "vlseg4e8[ff].v,e32,m4";
	    34'b0000111???????101?01001000?0000011  :  Instruction = "vlseg4e16[ff].v,e32,m4";
	    34'b0000111???????000?01001100?0000011  :  Instruction = "vlseg4e8[ff].v,e32,m8";
	    34'b0000111???????110?01010110?????011  :  Instruction = "vlsseg4e32.v,e32,mf8";
	    34'b0000111???????111?01010110?????011  :  Instruction = "vlsseg4e64.v,e32,mf8";
	    34'b0000111???????101?01011010?????011  :  Instruction = "vlsseg4e16.v,e32,mf4";
	    34'b0000111???????110?01011010?????011  :  Instruction = "vlsseg4e32.v,e32,mf4";
	    34'b0000111???????111?01011010?????011  :  Instruction = "vlsseg4e64.v,e32,mf4";
	    34'b0000111???????000?01011110?????011  :  Instruction = "vlsseg4e8.v,e32,mf2";
	    34'b0000111???????101?01011110?????011  :  Instruction = "vlsseg4e16.v,e32,mf2";
	    34'b0000111???????110?01011110?????011  :  Instruction = "vlsseg4e32.v,e32,mf2";
	    34'b0000111???????111?01011110?????011  :  Instruction = "vlsseg4e64.v,e32,mf2";
	    34'b0000111???????000?01000010?????011  :  Instruction = "vlsseg4e8.v,e32,m1";
	    34'b0000111???????101?01000010?????011  :  Instruction = "vlsseg4e16.v,e32,m1";
	    34'b0000111???????110?01000010?????011  :  Instruction = "vlsseg4e32.v,e32,m1";
	    34'b0000111???????111?01000010?????011  :  Instruction = "vlsseg4e64.v,e32,m1";
	    34'b0000111???????000?01000110?????011  :  Instruction = "vlsseg4e8.v,e32,m2";
	    34'b0000111???????101?01000110?????011  :  Instruction = "vlsseg4e16.v,e32,m2";
	    34'b0000111???????110?01000110?????011  :  Instruction = "vlsseg4e32.v,e32,m2";
	    34'b0000111???????000?01001010?????011  :  Instruction = "vlsseg4e8.v,e32,m4";
	    34'b0000111???????101?01001010?????011  :  Instruction = "vlsseg4e16.v,e32,m4";
	    34'b0000111???????000?01001110?????011  :  Instruction = "vlsseg4e8.v,e32,m8";
	    34'b0000111???????000?010???0001000011  :  Instruction = "vl4re8.v,e32";
	    34'b0000111???????101?010???0001000011  :  Instruction = "vl4re16.v,e32";
	    34'b0000111???????110?010???0001000011  :  Instruction = "vl4re32.v,e32";
	    34'b0000111???????111?010???0001000011  :  Instruction = "vl4re64.v,e32";
	    34'b0000111???????110?010101?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e32,mf8";
	    34'b0000111???????111?010101?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e32,mf8";
	    34'b0000111???????101?010110?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e32,mf4";
	    34'b0000111???????110?010110?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e32,mf4";
	    34'b0000111???????111?010110?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e32,mf4";
	    34'b0000111???????000?010111?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e32,mf2";
	    34'b0000111???????101?010111?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e32,mf2";
	    34'b0000111???????110?010111?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e32,mf2";
	    34'b0000111???????111?010111?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e32,mf2";
	    34'b0000111???????000?010000?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e32,m1";
	    34'b0000111???????101?010000?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e32,m1";
	    34'b0000111???????110?010000?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e32,m1";
	    34'b0000111???????111?010000?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e32,m1";
	    34'b0000111???????000?010001?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e32,m2";
	    34'b0000111???????101?010001?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e32,m2";
	    34'b0000111???????110?010001?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e32,m2";
	    34'b0000111???????111?010001?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e32,m2";
	    34'b0000111???????110?01010100?0000100  :  Instruction = "vlseg5e32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000100  :  Instruction = "vlseg5e64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000100  :  Instruction = "vlseg5e16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000100  :  Instruction = "vlseg5e32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000100  :  Instruction = "vlseg5e64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000100  :  Instruction = "vlseg5e8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000100  :  Instruction = "vlseg5e16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000100  :  Instruction = "vlseg5e32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000100  :  Instruction = "vlseg5e64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000100  :  Instruction = "vlseg5e8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000100  :  Instruction = "vlseg5e16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000100  :  Instruction = "vlseg5e32[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000100  :  Instruction = "vlseg5e8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000100  :  Instruction = "vlseg5e16[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000100  :  Instruction = "vlseg5e8[ff].v,e32,m4";
	    34'b0000111???????110?01010110?????100  :  Instruction = "vlsseg5e32.v,e32,mf8";
	    34'b0000111???????111?01010110?????100  :  Instruction = "vlsseg5e64.v,e32,mf8";
	    34'b0000111???????101?01011010?????100  :  Instruction = "vlsseg5e16.v,e32,mf4";
	    34'b0000111???????110?01011010?????100  :  Instruction = "vlsseg5e32.v,e32,mf4";
	    34'b0000111???????111?01011010?????100  :  Instruction = "vlsseg5e64.v,e32,mf4";
	    34'b0000111???????000?01011110?????100  :  Instruction = "vlsseg5e8.v,e32,mf2";
	    34'b0000111???????101?01011110?????100  :  Instruction = "vlsseg5e16.v,e32,mf2";
	    34'b0000111???????110?01011110?????100  :  Instruction = "vlsseg5e32.v,e32,mf2";
	    34'b0000111???????111?01011110?????100  :  Instruction = "vlsseg5e64.v,e32,mf2";
	    34'b0000111???????000?01000010?????100  :  Instruction = "vlsseg5e8.v,e32,m1";
	    34'b0000111???????101?01000010?????100  :  Instruction = "vlsseg5e16.v,e32,m1";
	    34'b0000111???????110?01000010?????100  :  Instruction = "vlsseg5e32.v,e32,m1";
	    34'b0000111???????000?01000110?????100  :  Instruction = "vlsseg5e8.v,e32,m2";
	    34'b0000111???????101?01000110?????100  :  Instruction = "vlsseg5e16.v,e32,m2";
	    34'b0000111???????000?01001010?????100  :  Instruction = "vlsseg5e8.v,e32,m4";
	    34'b0000111???????110?010101?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e32,mf8";
	    34'b0000111???????111?010101?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e32,mf8";
	    34'b0000111???????101?010110?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e32,mf4";
	    34'b0000111???????110?010110?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e32,mf4";
	    34'b0000111???????111?010110?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e32,mf4";
	    34'b0000111???????000?010111?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e32,mf2";
	    34'b0000111???????101?010111?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e32,mf2";
	    34'b0000111???????110?010111?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e32,mf2";
	    34'b0000111???????111?010111?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e32,mf2";
	    34'b0000111???????000?010000?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e32,m1";
	    34'b0000111???????101?010000?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e32,m1";
	    34'b0000111???????110?010000?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e32,m1";
	    34'b0000111???????111?010000?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e32,m1";
	    34'b0000111???????110?01010100?0000101  :  Instruction = "vlseg6e32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000101  :  Instruction = "vlseg6e64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000101  :  Instruction = "vlseg6e16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000101  :  Instruction = "vlseg6e32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000101  :  Instruction = "vlseg6e64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000101  :  Instruction = "vlseg6e8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000101  :  Instruction = "vlseg6e16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000101  :  Instruction = "vlseg6e32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000101  :  Instruction = "vlseg6e64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000101  :  Instruction = "vlseg6e8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000101  :  Instruction = "vlseg6e16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000101  :  Instruction = "vlseg6e32[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000101  :  Instruction = "vlseg6e8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000101  :  Instruction = "vlseg6e16[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000101  :  Instruction = "vlseg6e8[ff].v,e32,m4";
	    34'b0000111???????110?01010110?????101  :  Instruction = "vlsseg6e32.v,e32,mf8";
	    34'b0000111???????111?01010110?????101  :  Instruction = "vlsseg6e64.v,e32,mf8";
	    34'b0000111???????101?01011010?????101  :  Instruction = "vlsseg6e16.v,e32,mf4";
	    34'b0000111???????110?01011010?????101  :  Instruction = "vlsseg6e32.v,e32,mf4";
	    34'b0000111???????111?01011010?????101  :  Instruction = "vlsseg6e64.v,e32,mf4";
	    34'b0000111???????000?01011110?????101  :  Instruction = "vlsseg6e8.v,e32,mf2";
	    34'b0000111???????101?01011110?????101  :  Instruction = "vlsseg6e16.v,e32,mf2";
	    34'b0000111???????110?01011110?????101  :  Instruction = "vlsseg6e32.v,e32,mf2";
	    34'b0000111???????111?01011110?????101  :  Instruction = "vlsseg6e64.v,e32,mf2";
	    34'b0000111???????000?01000010?????101  :  Instruction = "vlsseg6e8.v,e32,m1";
	    34'b0000111???????101?01000010?????101  :  Instruction = "vlsseg6e16.v,e32,m1";
	    34'b0000111???????110?01000010?????101  :  Instruction = "vlsseg6e32.v,e32,m1";
	    34'b0000111???????000?01000110?????101  :  Instruction = "vlsseg6e8.v,e32,m2";
	    34'b0000111???????101?01000110?????101  :  Instruction = "vlsseg6e16.v,e32,m2";
	    34'b0000111???????000?01001010?????101  :  Instruction = "vlsseg6e8.v,e32,m4";
	    34'b0000111???????110?010101?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e32,mf8";
	    34'b0000111???????111?010101?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e32,mf8";
	    34'b0000111???????101?010110?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e32,mf4";
	    34'b0000111???????110?010110?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e32,mf4";
	    34'b0000111???????111?010110?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e32,mf4";
	    34'b0000111???????000?010111?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e32,mf2";
	    34'b0000111???????101?010111?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e32,mf2";
	    34'b0000111???????110?010111?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e32,mf2";
	    34'b0000111???????111?010111?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e32,mf2";
	    34'b0000111???????000?010000?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e32,m1";
	    34'b0000111???????101?010000?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e32,m1";
	    34'b0000111???????110?010000?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e32,m1";
	    34'b0000111???????111?010000?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e32,m1";
	    34'b0000111???????110?01010100?0000110  :  Instruction = "vlseg7e32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000110  :  Instruction = "vlseg7e64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000110  :  Instruction = "vlseg7e16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000110  :  Instruction = "vlseg7e32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000110  :  Instruction = "vlseg7e64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000110  :  Instruction = "vlseg7e8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000110  :  Instruction = "vlseg7e16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000110  :  Instruction = "vlseg7e32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000110  :  Instruction = "vlseg7e64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000110  :  Instruction = "vlseg7e8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000110  :  Instruction = "vlseg7e16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000110  :  Instruction = "vlseg7e32[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000110  :  Instruction = "vlseg7e8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000110  :  Instruction = "vlseg7e16[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000110  :  Instruction = "vlseg7e8[ff].v,e32,m4";
	    34'b0000111???????110?01010110?????110  :  Instruction = "vlsseg7e32.v,e32,mf8";
	    34'b0000111???????111?01010110?????110  :  Instruction = "vlsseg7e64.v,e32,mf8";
	    34'b0000111???????101?01011010?????110  :  Instruction = "vlsseg7e16.v,e32,mf4";
	    34'b0000111???????110?01011010?????110  :  Instruction = "vlsseg7e32.v,e32,mf4";
	    34'b0000111???????111?01011010?????110  :  Instruction = "vlsseg7e64.v,e32,mf4";
	    34'b0000111???????000?01011110?????110  :  Instruction = "vlsseg7e8.v,e32,mf2";
	    34'b0000111???????101?01011110?????110  :  Instruction = "vlsseg7e16.v,e32,mf2";
	    34'b0000111???????110?01011110?????110  :  Instruction = "vlsseg7e32.v,e32,mf2";
	    34'b0000111???????111?01011110?????110  :  Instruction = "vlsseg7e64.v,e32,mf2";
	    34'b0000111???????000?01000010?????110  :  Instruction = "vlsseg7e8.v,e32,m1";
	    34'b0000111???????101?01000010?????110  :  Instruction = "vlsseg7e16.v,e32,m1";
	    34'b0000111???????110?01000010?????110  :  Instruction = "vlsseg7e32.v,e32,m1";
	    34'b0000111???????000?01000110?????110  :  Instruction = "vlsseg7e8.v,e32,m2";
	    34'b0000111???????101?01000110?????110  :  Instruction = "vlsseg7e16.v,e32,m2";
	    34'b0000111???????000?01001010?????110  :  Instruction = "vlsseg7e8.v,e32,m4";
	    34'b0000111???????110?010101?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e32,mf8";
	    34'b0000111???????111?010101?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e32,mf8";
	    34'b0000111???????101?010110?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e32,mf4";
	    34'b0000111???????110?010110?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e32,mf4";
	    34'b0000111???????111?010110?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e32,mf4";
	    34'b0000111???????000?010111?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e32,mf2";
	    34'b0000111???????101?010111?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e32,mf2";
	    34'b0000111???????110?010111?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e32,mf2";
	    34'b0000111???????111?010111?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e32,mf2";
	    34'b0000111???????000?010000?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e32,m1";
	    34'b0000111???????101?010000?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e32,m1";
	    34'b0000111???????110?010000?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e32,m1";
	    34'b0000111???????111?010000?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e32,m1";
	    34'b0000111???????110?01010100?0000111  :  Instruction = "vlseg8e32[ff].v,e32,mf8";
	    34'b0000111???????111?01010100?0000111  :  Instruction = "vlseg8e64[ff].v,e32,mf8";
	    34'b0000111???????101?01011000?0000111  :  Instruction = "vlseg8e16[ff].v,e32,mf4";
	    34'b0000111???????110?01011000?0000111  :  Instruction = "vlseg8e32[ff].v,e32,mf4";
	    34'b0000111???????111?01011000?0000111  :  Instruction = "vlseg8e64[ff].v,e32,mf4";
	    34'b0000111???????000?01011100?0000111  :  Instruction = "vlseg8e8[ff].v,e32,mf2";
	    34'b0000111???????101?01011100?0000111  :  Instruction = "vlseg8e16[ff].v,e32,mf2";
	    34'b0000111???????110?01011100?0000111  :  Instruction = "vlseg8e32[ff].v,e32,mf2";
	    34'b0000111???????111?01011100?0000111  :  Instruction = "vlseg8e64[ff].v,e32,mf2";
	    34'b0000111???????000?01000000?0000111  :  Instruction = "vlseg8e8[ff].v,e32,m1";
	    34'b0000111???????101?01000000?0000111  :  Instruction = "vlseg8e16[ff].v,e32,m1";
	    34'b0000111???????110?01000000?0000111  :  Instruction = "vlseg8e32[ff].v,e32,m1";
	    34'b0000111???????000?01000100?0000111  :  Instruction = "vlseg8e8[ff].v,e32,m2";
	    34'b0000111???????101?01000100?0000111  :  Instruction = "vlseg8e16[ff].v,e32,m2";
	    34'b0000111???????000?01001000?0000111  :  Instruction = "vlseg8e8[ff].v,e32,m4";
	    34'b0000111???????000?010???0001000111  :  Instruction = "vl8re8.v,e32";
	    34'b0000111???????101?010???0001000111  :  Instruction = "vl8re16.v,e32";
	    34'b0000111???????110?010???0001000111  :  Instruction = "vl8re32.v,e32";
	    34'b0000111???????111?010???0001000111  :  Instruction = "vl8re64.v,e32";
	    34'b0000111???????110?01010110?????111  :  Instruction = "vlsseg8e32.v,e32,mf8";
	    34'b0000111???????111?01010110?????111  :  Instruction = "vlsseg8e64.v,e32,mf8";
	    34'b0000111???????101?01011010?????111  :  Instruction = "vlsseg8e16.v,e32,mf4";
	    34'b0000111???????110?01011010?????111  :  Instruction = "vlsseg8e32.v,e32,mf4";
	    34'b0000111???????111?01011010?????111  :  Instruction = "vlsseg8e64.v,e32,mf4";
	    34'b0000111???????000?01011110?????111  :  Instruction = "vlsseg8e8.v,e32,mf2";
	    34'b0000111???????101?01011110?????111  :  Instruction = "vlsseg8e16.v,e32,mf2";
	    34'b0000111???????110?01011110?????111  :  Instruction = "vlsseg8e32.v,e32,mf2";
	    34'b0000111???????111?01011110?????111  :  Instruction = "vlsseg8e64.v,e32,mf2";
	    34'b0000111???????000?01000010?????111  :  Instruction = "vlsseg8e8.v,e32,m1";
	    34'b0000111???????101?01000010?????111  :  Instruction = "vlsseg8e16.v,e32,m1";
	    34'b0000111???????110?01000010?????111  :  Instruction = "vlsseg8e32.v,e32,m1";
	    34'b0000111???????000?01000110?????111  :  Instruction = "vlsseg8e8.v,e32,m2";
	    34'b0000111???????101?01000110?????111  :  Instruction = "vlsseg8e16.v,e32,m2";
	    34'b0000111???????000?01001010?????111  :  Instruction = "vlsseg8e8.v,e32,m4";
	    34'b0000111???????110?010101?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e32,mf8";
	    34'b0000111???????111?010101?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e32,mf8";
	    34'b0000111???????101?010110?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e32,mf4";
	    34'b0000111???????110?010110?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e32,mf4";
	    34'b0000111???????111?010110?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e32,mf4";
	    34'b0000111???????000?010111?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e32,mf2";
	    34'b0000111???????101?010111?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e32,mf2";
	    34'b0000111???????110?010111?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e32,mf2";
	    34'b0000111???????111?010111?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e32,mf2";
	    34'b0000111???????000?010000?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e32,m1";
	    34'b0000111???????101?010000?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e32,m1";
	    34'b0000111???????110?010000?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e32,m1";
	    34'b0000111???????111?010000?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e32,m1";
	    34'b0100111???????110?01010100?0000???  :  Instruction = "vse32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000???  :  Instruction = "vse64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000???  :  Instruction = "vse16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000???  :  Instruction = "vse32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000???  :  Instruction = "vse64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000???  :  Instruction = "vse8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000???  :  Instruction = "vse16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000???  :  Instruction = "vse32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000???  :  Instruction = "vse64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000???  :  Instruction = "vse8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000???  :  Instruction = "vse16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000???  :  Instruction = "vse32[ff].v,e32,m1";
	    34'b0100111???????111?01000000?0000???  :  Instruction = "vse64[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000???  :  Instruction = "vse8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000???  :  Instruction = "vse16[ff].v,e32,m2";
	    34'b0100111???????110?01000100?0000???  :  Instruction = "vse32[ff].v,e32,m2";
	    34'b0100111???????111?01000100?0000???  :  Instruction = "vse64[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000???  :  Instruction = "vse8[ff].v,e32,m4";
	    34'b0100111???????101?01001000?0000???  :  Instruction = "vse16[ff].v,e32,m4";
	    34'b0100111???????110?01001000?0000???  :  Instruction = "vse32[ff].v,e32,m4";
	    34'b0100111???????111?01001000?0000???  :  Instruction = "vse64[ff].v,e32,m4";
	    34'b0100111???????000?01001100?0000???  :  Instruction = "vse8[ff].v,e32,m8";
	    34'b0100111???????101?01001100?0000???  :  Instruction = "vse16[ff].v,e32,m8";
	    34'b0100111???????110?01001100?0000???  :  Instruction = "vse32[ff].v,e32,m8";
	    34'b0100111???????000?010???0001000000  :  Instruction = "vs1r.v,e32";
	    34'b0100111???????110?01010110????????  :  Instruction = "vsse32.v,e32,mf8";
	    34'b0100111???????111?01010110????????  :  Instruction = "vsse64.v,e32,mf8";
	    34'b0100111???????101?01011010????????  :  Instruction = "vsse16.v,e32,mf4";
	    34'b0100111???????110?01011010????????  :  Instruction = "vsse32.v,e32,mf4";
	    34'b0100111???????111?01011010????????  :  Instruction = "vsse64.v,e32,mf4";
	    34'b0100111???????000?01011110????????  :  Instruction = "vsse8.v,e32,mf2";
	    34'b0100111???????101?01011110????????  :  Instruction = "vsse16.v,e32,mf2";
	    34'b0100111???????110?01011110????????  :  Instruction = "vsse32.v,e32,mf2";
	    34'b0100111???????111?01011110????????  :  Instruction = "vsse64.v,e32,mf2";
	    34'b0100111???????000?01000010????????  :  Instruction = "vsse8.v,e32,m1";
	    34'b0100111???????101?01000010????????  :  Instruction = "vsse16.v,e32,m1";
	    34'b0100111???????110?01000010????????  :  Instruction = "vsse32.v,e32,m1";
	    34'b0100111???????111?01000010????????  :  Instruction = "vsse64.v,e32,m1";
	    34'b0100111???????000?01000110????????  :  Instruction = "vsse8.v,e32,m2";
	    34'b0100111???????101?01000110????????  :  Instruction = "vsse16.v,e32,m2";
	    34'b0100111???????110?01000110????????  :  Instruction = "vsse32.v,e32,m2";
	    34'b0100111???????111?01000110????????  :  Instruction = "vsse64.v,e32,m2";
	    34'b0100111???????000?01001010????????  :  Instruction = "vsse8.v,e32,m4";
	    34'b0100111???????101?01001010????????  :  Instruction = "vsse16.v,e32,m4";
	    34'b0100111???????110?01001010????????  :  Instruction = "vsse32.v,e32,m4";
	    34'b0100111???????111?01001010????????  :  Instruction = "vsse64.v,e32,m4";
	    34'b0100111???????000?01001110????????  :  Instruction = "vsse8.v,e32,m8";
	    34'b0100111???????101?01001110????????  :  Instruction = "vsse16.v,e32,m8";
	    34'b0100111???????110?01001110????????  :  Instruction = "vsse32.v,e32,m8";
	    34'b0100111???????110?010101?1????????  :  Instruction = "vs[uo]xei32.v,e32,mf8";
	    34'b0100111???????111?010101?1????????  :  Instruction = "vs[uo]xei64.v,e32,mf8";
	    34'b0100111???????101?010110?1????????  :  Instruction = "vs[uo]xei16.v,e32,mf4";
	    34'b0100111???????110?010110?1????????  :  Instruction = "vs[uo]xei32.v,e32,mf4";
	    34'b0100111???????111?010110?1????????  :  Instruction = "vs[uo]xei64.v,e32,mf4";
	    34'b0100111???????000?010111?1????????  :  Instruction = "vs[uo]xei8.v,e32,mf2";
	    34'b0100111???????101?010111?1????????  :  Instruction = "vs[uo]xei16.v,e32,mf2";
	    34'b0100111???????110?010111?1????????  :  Instruction = "vs[uo]xei32.v,e32,mf2";
	    34'b0100111???????111?010111?1????????  :  Instruction = "vs[uo]xei64.v,e32,mf2";
	    34'b0100111???????000?010000?1????????  :  Instruction = "vs[uo]xei8.v,e32,m1";
	    34'b0100111???????101?010000?1????????  :  Instruction = "vs[uo]xei16.v,e32,m1";
	    34'b0100111???????110?010000?1????????  :  Instruction = "vs[uo]xei32.v,e32,m1";
	    34'b0100111???????111?010000?1????????  :  Instruction = "vs[uo]xei64.v,e32,m1";
	    34'b0100111???????000?010001?1????????  :  Instruction = "vs[uo]xei8.v,e32,m2";
	    34'b0100111???????101?010001?1????????  :  Instruction = "vs[uo]xei16.v,e32,m2";
	    34'b0100111???????110?010001?1????????  :  Instruction = "vs[uo]xei32.v,e32,m2";
	    34'b0100111???????111?010001?1????????  :  Instruction = "vs[uo]xei64.v,e32,m2";
	    34'b0100111???????000?010010?1????????  :  Instruction = "vs[uo]xei8.v,e32,m4";
	    34'b0100111???????101?010010?1????????  :  Instruction = "vs[uo]xei16.v,e32,m4";
	    34'b0100111???????110?010010?1????????  :  Instruction = "vs[uo]xei32.v,e32,m4";
	    34'b0100111???????111?010010?1????????  :  Instruction = "vs[uo]xei64.v,e32,m4";
	    34'b0100111???????000?010011?1????????  :  Instruction = "vs[uo]xei8.v,e32,m8";
	    34'b0100111???????101?010011?1????????  :  Instruction = "vs[uo]xei16.v,e32,m8";
	    34'b0100111???????110?010011?1????????  :  Instruction = "vs[uo]xei32.v,e32,m8";
	    34'b0100111???????110?01010100?0000001  :  Instruction = "vsseg2e32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000001  :  Instruction = "vsseg2e64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000001  :  Instruction = "vsseg2e16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000001  :  Instruction = "vsseg2e32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000001  :  Instruction = "vsseg2e64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000001  :  Instruction = "vsseg2e8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000001  :  Instruction = "vsseg2e16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000001  :  Instruction = "vsseg2e32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000001  :  Instruction = "vsseg2e64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000001  :  Instruction = "vsseg2e8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000001  :  Instruction = "vsseg2e16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000001  :  Instruction = "vsseg2e32[ff].v,e32,m1";
	    34'b0100111???????111?01000000?0000001  :  Instruction = "vsseg2e64[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000001  :  Instruction = "vsseg2e8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000001  :  Instruction = "vsseg2e16[ff].v,e32,m2";
	    34'b0100111???????110?01000100?0000001  :  Instruction = "vsseg2e32[ff].v,e32,m2";
	    34'b0100111???????111?01000100?0000001  :  Instruction = "vsseg2e64[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000001  :  Instruction = "vsseg2e8[ff].v,e32,m4";
	    34'b0100111???????101?01001000?0000001  :  Instruction = "vsseg2e16[ff].v,e32,m4";
	    34'b0100111???????110?01001000?0000001  :  Instruction = "vsseg2e32[ff].v,e32,m4";
	    34'b0100111???????000?01001100?0000001  :  Instruction = "vsseg2e8[ff].v,e32,m8";
	    34'b0100111???????101?01001100?0000001  :  Instruction = "vsseg2e16[ff].v,e32,m8";
	    34'b0100111???????000?010???0001000001  :  Instruction = "vs2r.v,e32";
	    34'b0100111???????110?01010110?????001  :  Instruction = "vssseg2e32.v,e32,mf8";
	    34'b0100111???????111?01010110?????001  :  Instruction = "vssseg2e64.v,e32,mf8";
	    34'b0100111???????101?01011010?????001  :  Instruction = "vssseg2e16.v,e32,mf4";
	    34'b0100111???????110?01011010?????001  :  Instruction = "vssseg2e32.v,e32,mf4";
	    34'b0100111???????111?01011010?????001  :  Instruction = "vssseg2e64.v,e32,mf4";
	    34'b0100111???????000?01011110?????001  :  Instruction = "vssseg2e8.v,e32,mf2";
	    34'b0100111???????101?01011110?????001  :  Instruction = "vssseg2e16.v,e32,mf2";
	    34'b0100111???????110?01011110?????001  :  Instruction = "vssseg2e32.v,e32,mf2";
	    34'b0100111???????111?01011110?????001  :  Instruction = "vssseg2e64.v,e32,mf2";
	    34'b0100111???????000?01000010?????001  :  Instruction = "vssseg2e8.v,e32,m1";
	    34'b0100111???????101?01000010?????001  :  Instruction = "vssseg2e16.v,e32,m1";
	    34'b0100111???????110?01000010?????001  :  Instruction = "vssseg2e32.v,e32,m1";
	    34'b0100111???????111?01000010?????001  :  Instruction = "vssseg2e64.v,e32,m1";
	    34'b0100111???????000?01000110?????001  :  Instruction = "vssseg2e8.v,e32,m2";
	    34'b0100111???????101?01000110?????001  :  Instruction = "vssseg2e16.v,e32,m2";
	    34'b0100111???????110?01000110?????001  :  Instruction = "vssseg2e32.v,e32,m2";
	    34'b0100111???????111?01000110?????001  :  Instruction = "vssseg2e64.v,e32,m2";
	    34'b0100111???????000?01001010?????001  :  Instruction = "vssseg2e8.v,e32,m4";
	    34'b0100111???????101?01001010?????001  :  Instruction = "vssseg2e16.v,e32,m4";
	    34'b0100111???????110?01001010?????001  :  Instruction = "vssseg2e32.v,e32,m4";
	    34'b0100111???????000?01001110?????001  :  Instruction = "vssseg2e8.v,e32,m8";
	    34'b0100111???????101?01001110?????001  :  Instruction = "vssseg2e16.v,e32,m8";
	    34'b0100111???????110?010101?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e32,mf8";
	    34'b0100111???????111?010101?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e32,mf8";
	    34'b0100111???????101?010110?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e32,mf4";
	    34'b0100111???????110?010110?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e32,mf4";
	    34'b0100111???????111?010110?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e32,mf4";
	    34'b0100111???????000?010111?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e32,mf2";
	    34'b0100111???????101?010111?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e32,mf2";
	    34'b0100111???????110?010111?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e32,mf2";
	    34'b0100111???????111?010111?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e32,mf2";
	    34'b0100111???????000?010000?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e32,m1";
	    34'b0100111???????101?010000?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e32,m1";
	    34'b0100111???????110?010000?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e32,m1";
	    34'b0100111???????111?010000?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e32,m1";
	    34'b0100111???????000?010001?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e32,m2";
	    34'b0100111???????101?010001?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e32,m2";
	    34'b0100111???????110?010001?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e32,m2";
	    34'b0100111???????111?010001?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e32,m2";
	    34'b0100111???????000?010010?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e32,m4";
	    34'b0100111???????101?010010?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e32,m4";
	    34'b0100111???????110?010010?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e32,m4";
	    34'b0100111???????111?010010?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e32,m4";
	    34'b0100111???????110?01010100?0000010  :  Instruction = "vsseg3e32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000010  :  Instruction = "vsseg3e64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000010  :  Instruction = "vsseg3e16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000010  :  Instruction = "vsseg3e32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000010  :  Instruction = "vsseg3e64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000010  :  Instruction = "vsseg3e8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000010  :  Instruction = "vsseg3e16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000010  :  Instruction = "vsseg3e32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000010  :  Instruction = "vsseg3e64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000010  :  Instruction = "vsseg3e8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000010  :  Instruction = "vsseg3e16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000010  :  Instruction = "vsseg3e32[ff].v,e32,m1";
	    34'b0100111???????111?01000000?0000010  :  Instruction = "vsseg3e64[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000010  :  Instruction = "vsseg3e8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000010  :  Instruction = "vsseg3e16[ff].v,e32,m2";
	    34'b0100111???????110?01000100?0000010  :  Instruction = "vsseg3e32[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000010  :  Instruction = "vsseg3e8[ff].v,e32,m4";
	    34'b0100111???????101?01001000?0000010  :  Instruction = "vsseg3e16[ff].v,e32,m4";
	    34'b0100111???????000?01001100?0000010  :  Instruction = "vsseg3e8[ff].v,e32,m8";
	    34'b0100111???????110?01010110?????010  :  Instruction = "vssseg3e32.v,e32,mf8";
	    34'b0100111???????111?01010110?????010  :  Instruction = "vssseg3e64.v,e32,mf8";
	    34'b0100111???????101?01011010?????010  :  Instruction = "vssseg3e16.v,e32,mf4";
	    34'b0100111???????110?01011010?????010  :  Instruction = "vssseg3e32.v,e32,mf4";
	    34'b0100111???????111?01011010?????010  :  Instruction = "vssseg3e64.v,e32,mf4";
	    34'b0100111???????000?01011110?????010  :  Instruction = "vssseg3e8.v,e32,mf2";
	    34'b0100111???????101?01011110?????010  :  Instruction = "vssseg3e16.v,e32,mf2";
	    34'b0100111???????110?01011110?????010  :  Instruction = "vssseg3e32.v,e32,mf2";
	    34'b0100111???????111?01011110?????010  :  Instruction = "vssseg3e64.v,e32,mf2";
	    34'b0100111???????000?01000010?????010  :  Instruction = "vssseg3e8.v,e32,m1";
	    34'b0100111???????101?01000010?????010  :  Instruction = "vssseg3e16.v,e32,m1";
	    34'b0100111???????110?01000010?????010  :  Instruction = "vssseg3e32.v,e32,m1";
	    34'b0100111???????111?01000010?????010  :  Instruction = "vssseg3e64.v,e32,m1";
	    34'b0100111???????000?01000110?????010  :  Instruction = "vssseg3e8.v,e32,m2";
	    34'b0100111???????101?01000110?????010  :  Instruction = "vssseg3e16.v,e32,m2";
	    34'b0100111???????110?01000110?????010  :  Instruction = "vssseg3e32.v,e32,m2";
	    34'b0100111???????000?01001010?????010  :  Instruction = "vssseg3e8.v,e32,m4";
	    34'b0100111???????101?01001010?????010  :  Instruction = "vssseg3e16.v,e32,m4";
	    34'b0100111???????000?01001110?????010  :  Instruction = "vssseg3e8.v,e32,m8";
	    34'b0100111???????110?010101?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e32,mf8";
	    34'b0100111???????111?010101?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e32,mf8";
	    34'b0100111???????101?010110?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e32,mf4";
	    34'b0100111???????110?010110?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e32,mf4";
	    34'b0100111???????111?010110?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e32,mf4";
	    34'b0100111???????000?010111?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e32,mf2";
	    34'b0100111???????101?010111?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e32,mf2";
	    34'b0100111???????110?010111?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e32,mf2";
	    34'b0100111???????111?010111?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e32,mf2";
	    34'b0100111???????000?010000?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e32,m1";
	    34'b0100111???????101?010000?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e32,m1";
	    34'b0100111???????110?010000?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e32,m1";
	    34'b0100111???????111?010000?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e32,m1";
	    34'b0100111???????000?010001?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e32,m2";
	    34'b0100111???????101?010001?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e32,m2";
	    34'b0100111???????110?010001?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e32,m2";
	    34'b0100111???????111?010001?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e32,m2";
	    34'b0100111???????110?01010100?0000011  :  Instruction = "vsseg4e32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000011  :  Instruction = "vsseg4e64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000011  :  Instruction = "vsseg4e16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000011  :  Instruction = "vsseg4e32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000011  :  Instruction = "vsseg4e64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000011  :  Instruction = "vsseg4e8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000011  :  Instruction = "vsseg4e16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000011  :  Instruction = "vsseg4e32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000011  :  Instruction = "vsseg4e64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000011  :  Instruction = "vsseg4e8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000011  :  Instruction = "vsseg4e16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000011  :  Instruction = "vsseg4e32[ff].v,e32,m1";
	    34'b0100111???????111?01000000?0000011  :  Instruction = "vsseg4e64[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000011  :  Instruction = "vsseg4e8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000011  :  Instruction = "vsseg4e16[ff].v,e32,m2";
	    34'b0100111???????110?01000100?0000011  :  Instruction = "vsseg4e32[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000011  :  Instruction = "vsseg4e8[ff].v,e32,m4";
	    34'b0100111???????101?01001000?0000011  :  Instruction = "vsseg4e16[ff].v,e32,m4";
	    34'b0100111???????000?01001100?0000011  :  Instruction = "vsseg4e8[ff].v,e32,m8";
	    34'b0100111???????110?01010110?????011  :  Instruction = "vssseg4e32.v,e32,mf8";
	    34'b0100111???????111?01010110?????011  :  Instruction = "vssseg4e64.v,e32,mf8";
	    34'b0100111???????101?01011010?????011  :  Instruction = "vssseg4e16.v,e32,mf4";
	    34'b0100111???????110?01011010?????011  :  Instruction = "vssseg4e32.v,e32,mf4";
	    34'b0100111???????111?01011010?????011  :  Instruction = "vssseg4e64.v,e32,mf4";
	    34'b0100111???????000?01011110?????011  :  Instruction = "vssseg4e8.v,e32,mf2";
	    34'b0100111???????101?01011110?????011  :  Instruction = "vssseg4e16.v,e32,mf2";
	    34'b0100111???????110?01011110?????011  :  Instruction = "vssseg4e32.v,e32,mf2";
	    34'b0100111???????111?01011110?????011  :  Instruction = "vssseg4e64.v,e32,mf2";
	    34'b0100111???????000?01000010?????011  :  Instruction = "vssseg4e8.v,e32,m1";
	    34'b0100111???????101?01000010?????011  :  Instruction = "vssseg4e16.v,e32,m1";
	    34'b0100111???????110?01000010?????011  :  Instruction = "vssseg4e32.v,e32,m1";
	    34'b0100111???????111?01000010?????011  :  Instruction = "vssseg4e64.v,e32,m1";
	    34'b0100111???????000?01000110?????011  :  Instruction = "vssseg4e8.v,e32,m2";
	    34'b0100111???????101?01000110?????011  :  Instruction = "vssseg4e16.v,e32,m2";
	    34'b0100111???????110?01000110?????011  :  Instruction = "vssseg4e32.v,e32,m2";
	    34'b0100111???????000?01001010?????011  :  Instruction = "vssseg4e8.v,e32,m4";
	    34'b0100111???????101?01001010?????011  :  Instruction = "vssseg4e16.v,e32,m4";
	    34'b0100111???????000?01001110?????011  :  Instruction = "vssseg4e8.v,e32,m8";
	    34'b0100111???????000?010???0001000011  :  Instruction = "vs4r.v,e32";
	    34'b0100111???????110?010101?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e32,mf8";
	    34'b0100111???????111?010101?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e32,mf8";
	    34'b0100111???????101?010110?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e32,mf4";
	    34'b0100111???????110?010110?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e32,mf4";
	    34'b0100111???????111?010110?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e32,mf4";
	    34'b0100111???????000?010111?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e32,mf2";
	    34'b0100111???????101?010111?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e32,mf2";
	    34'b0100111???????110?010111?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e32,mf2";
	    34'b0100111???????111?010111?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e32,mf2";
	    34'b0100111???????000?010000?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e32,m1";
	    34'b0100111???????101?010000?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e32,m1";
	    34'b0100111???????110?010000?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e32,m1";
	    34'b0100111???????111?010000?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e32,m1";
	    34'b0100111???????000?010001?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e32,m2";
	    34'b0100111???????101?010001?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e32,m2";
	    34'b0100111???????110?010001?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e32,m2";
	    34'b0100111???????111?010001?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e32,m2";
	    34'b0100111???????110?01010100?0000100  :  Instruction = "vsseg5e32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000100  :  Instruction = "vsseg5e64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000100  :  Instruction = "vsseg5e16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000100  :  Instruction = "vsseg5e32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000100  :  Instruction = "vsseg5e64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000100  :  Instruction = "vsseg5e8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000100  :  Instruction = "vsseg5e16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000100  :  Instruction = "vsseg5e32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000100  :  Instruction = "vsseg5e64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000100  :  Instruction = "vsseg5e8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000100  :  Instruction = "vsseg5e16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000100  :  Instruction = "vsseg5e32[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000100  :  Instruction = "vsseg5e8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000100  :  Instruction = "vsseg5e16[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000100  :  Instruction = "vsseg5e8[ff].v,e32,m4";
	    34'b0100111???????110?01010110?????100  :  Instruction = "vssseg5e32.v,e32,mf8";
	    34'b0100111???????111?01010110?????100  :  Instruction = "vssseg5e64.v,e32,mf8";
	    34'b0100111???????101?01011010?????100  :  Instruction = "vssseg5e16.v,e32,mf4";
	    34'b0100111???????110?01011010?????100  :  Instruction = "vssseg5e32.v,e32,mf4";
	    34'b0100111???????111?01011010?????100  :  Instruction = "vssseg5e64.v,e32,mf4";
	    34'b0100111???????000?01011110?????100  :  Instruction = "vssseg5e8.v,e32,mf2";
	    34'b0100111???????101?01011110?????100  :  Instruction = "vssseg5e16.v,e32,mf2";
	    34'b0100111???????110?01011110?????100  :  Instruction = "vssseg5e32.v,e32,mf2";
	    34'b0100111???????111?01011110?????100  :  Instruction = "vssseg5e64.v,e32,mf2";
	    34'b0100111???????000?01000010?????100  :  Instruction = "vssseg5e8.v,e32,m1";
	    34'b0100111???????101?01000010?????100  :  Instruction = "vssseg5e16.v,e32,m1";
	    34'b0100111???????110?01000010?????100  :  Instruction = "vssseg5e32.v,e32,m1";
	    34'b0100111???????000?01000110?????100  :  Instruction = "vssseg5e8.v,e32,m2";
	    34'b0100111???????101?01000110?????100  :  Instruction = "vssseg5e16.v,e32,m2";
	    34'b0100111???????000?01001010?????100  :  Instruction = "vssseg5e8.v,e32,m4";
	    34'b0100111???????110?010101?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e32,mf8";
	    34'b0100111???????111?010101?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e32,mf8";
	    34'b0100111???????101?010110?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e32,mf4";
	    34'b0100111???????110?010110?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e32,mf4";
	    34'b0100111???????111?010110?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e32,mf4";
	    34'b0100111???????000?010111?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e32,mf2";
	    34'b0100111???????101?010111?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e32,mf2";
	    34'b0100111???????110?010111?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e32,mf2";
	    34'b0100111???????111?010111?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e32,mf2";
	    34'b0100111???????000?010000?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e32,m1";
	    34'b0100111???????101?010000?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e32,m1";
	    34'b0100111???????110?010000?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e32,m1";
	    34'b0100111???????111?010000?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e32,m1";
	    34'b0100111???????110?01010100?0000101  :  Instruction = "vsseg6e32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000101  :  Instruction = "vsseg6e64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000101  :  Instruction = "vsseg6e16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000101  :  Instruction = "vsseg6e32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000101  :  Instruction = "vsseg6e64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000101  :  Instruction = "vsseg6e8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000101  :  Instruction = "vsseg6e16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000101  :  Instruction = "vsseg6e32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000101  :  Instruction = "vsseg6e64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000101  :  Instruction = "vsseg6e8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000101  :  Instruction = "vsseg6e16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000101  :  Instruction = "vsseg6e32[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000101  :  Instruction = "vsseg6e8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000101  :  Instruction = "vsseg6e16[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000101  :  Instruction = "vsseg6e8[ff].v,e32,m4";
	    34'b0100111???????110?01010110?????101  :  Instruction = "vssseg6e32.v,e32,mf8";
	    34'b0100111???????111?01010110?????101  :  Instruction = "vssseg6e64.v,e32,mf8";
	    34'b0100111???????101?01011010?????101  :  Instruction = "vssseg6e16.v,e32,mf4";
	    34'b0100111???????110?01011010?????101  :  Instruction = "vssseg6e32.v,e32,mf4";
	    34'b0100111???????111?01011010?????101  :  Instruction = "vssseg6e64.v,e32,mf4";
	    34'b0100111???????000?01011110?????101  :  Instruction = "vssseg6e8.v,e32,mf2";
	    34'b0100111???????101?01011110?????101  :  Instruction = "vssseg6e16.v,e32,mf2";
	    34'b0100111???????110?01011110?????101  :  Instruction = "vssseg6e32.v,e32,mf2";
	    34'b0100111???????111?01011110?????101  :  Instruction = "vssseg6e64.v,e32,mf2";
	    34'b0100111???????000?01000010?????101  :  Instruction = "vssseg6e8.v,e32,m1";
	    34'b0100111???????101?01000010?????101  :  Instruction = "vssseg6e16.v,e32,m1";
	    34'b0100111???????110?01000010?????101  :  Instruction = "vssseg6e32.v,e32,m1";
	    34'b0100111???????000?01000110?????101  :  Instruction = "vssseg6e8.v,e32,m2";
	    34'b0100111???????101?01000110?????101  :  Instruction = "vssseg6e16.v,e32,m2";
	    34'b0100111???????000?01001010?????101  :  Instruction = "vssseg6e8.v,e32,m4";
	    34'b0100111???????110?010101?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e32,mf8";
	    34'b0100111???????111?010101?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e32,mf8";
	    34'b0100111???????101?010110?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e32,mf4";
	    34'b0100111???????110?010110?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e32,mf4";
	    34'b0100111???????111?010110?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e32,mf4";
	    34'b0100111???????000?010111?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e32,mf2";
	    34'b0100111???????101?010111?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e32,mf2";
	    34'b0100111???????110?010111?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e32,mf2";
	    34'b0100111???????111?010111?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e32,mf2";
	    34'b0100111???????000?010000?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e32,m1";
	    34'b0100111???????101?010000?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e32,m1";
	    34'b0100111???????110?010000?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e32,m1";
	    34'b0100111???????111?010000?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e32,m1";
	    34'b0100111???????110?01010100?0000110  :  Instruction = "vsseg7e32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000110  :  Instruction = "vsseg7e64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000110  :  Instruction = "vsseg7e16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000110  :  Instruction = "vsseg7e32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000110  :  Instruction = "vsseg7e64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000110  :  Instruction = "vsseg7e8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000110  :  Instruction = "vsseg7e16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000110  :  Instruction = "vsseg7e32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000110  :  Instruction = "vsseg7e64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000110  :  Instruction = "vsseg7e8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000110  :  Instruction = "vsseg7e16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000110  :  Instruction = "vsseg7e32[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000110  :  Instruction = "vsseg7e8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000110  :  Instruction = "vsseg7e16[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000110  :  Instruction = "vsseg7e8[ff].v,e32,m4";
	    34'b0100111???????110?01010110?????110  :  Instruction = "vssseg7e32.v,e32,mf8";
	    34'b0100111???????111?01010110?????110  :  Instruction = "vssseg7e64.v,e32,mf8";
	    34'b0100111???????101?01011010?????110  :  Instruction = "vssseg7e16.v,e32,mf4";
	    34'b0100111???????110?01011010?????110  :  Instruction = "vssseg7e32.v,e32,mf4";
	    34'b0100111???????111?01011010?????110  :  Instruction = "vssseg7e64.v,e32,mf4";
	    34'b0100111???????000?01011110?????110  :  Instruction = "vssseg7e8.v,e32,mf2";
	    34'b0100111???????101?01011110?????110  :  Instruction = "vssseg7e16.v,e32,mf2";
	    34'b0100111???????110?01011110?????110  :  Instruction = "vssseg7e32.v,e32,mf2";
	    34'b0100111???????111?01011110?????110  :  Instruction = "vssseg7e64.v,e32,mf2";
	    34'b0100111???????000?01000010?????110  :  Instruction = "vssseg7e8.v,e32,m1";
	    34'b0100111???????101?01000010?????110  :  Instruction = "vssseg7e16.v,e32,m1";
	    34'b0100111???????110?01000010?????110  :  Instruction = "vssseg7e32.v,e32,m1";
	    34'b0100111???????000?01000110?????110  :  Instruction = "vssseg7e8.v,e32,m2";
	    34'b0100111???????101?01000110?????110  :  Instruction = "vssseg7e16.v,e32,m2";
	    34'b0100111???????000?01001010?????110  :  Instruction = "vssseg7e8.v,e32,m4";
	    34'b0100111???????110?010101?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e32,mf8";
	    34'b0100111???????111?010101?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e32,mf8";
	    34'b0100111???????101?010110?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e32,mf4";
	    34'b0100111???????110?010110?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e32,mf4";
	    34'b0100111???????111?010110?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e32,mf4";
	    34'b0100111???????000?010111?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e32,mf2";
	    34'b0100111???????101?010111?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e32,mf2";
	    34'b0100111???????110?010111?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e32,mf2";
	    34'b0100111???????111?010111?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e32,mf2";
	    34'b0100111???????000?010000?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e32,m1";
	    34'b0100111???????101?010000?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e32,m1";
	    34'b0100111???????110?010000?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e32,m1";
	    34'b0100111???????111?010000?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e32,m1";
	    34'b0100111???????110?01010100?0000111  :  Instruction = "vsseg8e32[ff].v,e32,mf8";
	    34'b0100111???????111?01010100?0000111  :  Instruction = "vsseg8e64[ff].v,e32,mf8";
	    34'b0100111???????101?01011000?0000111  :  Instruction = "vsseg8e16[ff].v,e32,mf4";
	    34'b0100111???????110?01011000?0000111  :  Instruction = "vsseg8e32[ff].v,e32,mf4";
	    34'b0100111???????111?01011000?0000111  :  Instruction = "vsseg8e64[ff].v,e32,mf4";
	    34'b0100111???????000?01011100?0000111  :  Instruction = "vsseg8e8[ff].v,e32,mf2";
	    34'b0100111???????101?01011100?0000111  :  Instruction = "vsseg8e16[ff].v,e32,mf2";
	    34'b0100111???????110?01011100?0000111  :  Instruction = "vsseg8e32[ff].v,e32,mf2";
	    34'b0100111???????111?01011100?0000111  :  Instruction = "vsseg8e64[ff].v,e32,mf2";
	    34'b0100111???????000?01000000?0000111  :  Instruction = "vsseg8e8[ff].v,e32,m1";
	    34'b0100111???????101?01000000?0000111  :  Instruction = "vsseg8e16[ff].v,e32,m1";
	    34'b0100111???????110?01000000?0000111  :  Instruction = "vsseg8e32[ff].v,e32,m1";
	    34'b0100111???????000?01000100?0000111  :  Instruction = "vsseg8e8[ff].v,e32,m2";
	    34'b0100111???????101?01000100?0000111  :  Instruction = "vsseg8e16[ff].v,e32,m2";
	    34'b0100111???????000?01001000?0000111  :  Instruction = "vsseg8e8[ff].v,e32,m4";
	    34'b0100111???????000?010???0001000111  :  Instruction = "vs8r.v,e32";
	    34'b0100111???????110?01010110?????111  :  Instruction = "vssseg8e32.v,e32,mf8";
	    34'b0100111???????111?01010110?????111  :  Instruction = "vssseg8e64.v,e32,mf8";
	    34'b0100111???????101?01011010?????111  :  Instruction = "vssseg8e16.v,e32,mf4";
	    34'b0100111???????110?01011010?????111  :  Instruction = "vssseg8e32.v,e32,mf4";
	    34'b0100111???????111?01011010?????111  :  Instruction = "vssseg8e64.v,e32,mf4";
	    34'b0100111???????000?01011110?????111  :  Instruction = "vssseg8e8.v,e32,mf2";
	    34'b0100111???????101?01011110?????111  :  Instruction = "vssseg8e16.v,e32,mf2";
	    34'b0100111???????110?01011110?????111  :  Instruction = "vssseg8e32.v,e32,mf2";
	    34'b0100111???????111?01011110?????111  :  Instruction = "vssseg8e64.v,e32,mf2";
	    34'b0100111???????000?01000010?????111  :  Instruction = "vssseg8e8.v,e32,m1";
	    34'b0100111???????101?01000010?????111  :  Instruction = "vssseg8e16.v,e32,m1";
	    34'b0100111???????110?01000010?????111  :  Instruction = "vssseg8e32.v,e32,m1";
	    34'b0100111???????000?01000110?????111  :  Instruction = "vssseg8e8.v,e32,m2";
	    34'b0100111???????101?01000110?????111  :  Instruction = "vssseg8e16.v,e32,m2";
	    34'b0100111???????000?01001010?????111  :  Instruction = "vssseg8e8.v,e32,m4";
	    34'b0100111???????110?010101?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e32,mf8";
	    34'b0100111???????111?010101?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e32,mf8";
	    34'b0100111???????101?010110?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e32,mf4";
	    34'b0100111???????110?010110?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e32,mf4";
	    34'b0100111???????111?010110?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e32,mf4";
	    34'b0100111???????000?010111?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e32,mf2";
	    34'b0100111???????101?010111?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e32,mf2";
	    34'b0100111???????110?010111?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e32,mf2";
	    34'b0100111???????111?010111?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e32,mf2";
	    34'b0100111???????000?010000?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e32,m1";
	    34'b0100111???????101?010000?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e32,m1";
	    34'b0100111???????110?010000?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e32,m1";
	    34'b0100111???????111?010000?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e32,m1";
	    34'b0000111???????111?01110100?0000???  :  Instruction = "vle64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000???  :  Instruction = "vle32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000???  :  Instruction = "vle64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000???  :  Instruction = "vle16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000???  :  Instruction = "vle32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000???  :  Instruction = "vle64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000???  :  Instruction = "vle8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000???  :  Instruction = "vle16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000???  :  Instruction = "vle32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000???  :  Instruction = "vle64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000???  :  Instruction = "vle8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000???  :  Instruction = "vle16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000???  :  Instruction = "vle32[ff].v,e64,m2";
	    34'b0000111???????111?01100100?0000???  :  Instruction = "vle64[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000???  :  Instruction = "vle8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000???  :  Instruction = "vle16[ff].v,e64,m4";
	    34'b0000111???????110?01101000?0000???  :  Instruction = "vle32[ff].v,e64,m4";
	    34'b0000111???????111?01101000?0000???  :  Instruction = "vle64[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000???  :  Instruction = "vle8[ff].v,e64,m8";
	    34'b0000111???????101?01101100?0000???  :  Instruction = "vle16[ff].v,e64,m8";
	    34'b0000111???????110?01101100?0000???  :  Instruction = "vle32[ff].v,e64,m8";
	    34'b0000111???????111?01101100?0000???  :  Instruction = "vle64[ff].v,e64,m8";
	    34'b0000111???????000?011???0001000000  :  Instruction = "vl1re8.v,e64";
	    34'b0000111???????101?011???0001000000  :  Instruction = "vl1re16.v,e64";
	    34'b0000111???????110?011???0001000000  :  Instruction = "vl1re32.v,e64";
	    34'b0000111???????111?011???0001000000  :  Instruction = "vl1re64.v,e64";
	    34'b0000111???????111?01110110????????  :  Instruction = "vlse64.v,e64,mf8";
	    34'b0000111???????110?01111010????????  :  Instruction = "vlse32.v,e64,mf4";
	    34'b0000111???????111?01111010????????  :  Instruction = "vlse64.v,e64,mf4";
	    34'b0000111???????101?01111110????????  :  Instruction = "vlse16.v,e64,mf2";
	    34'b0000111???????110?01111110????????  :  Instruction = "vlse32.v,e64,mf2";
	    34'b0000111???????111?01111110????????  :  Instruction = "vlse64.v,e64,mf2";
	    34'b0000111???????000?01100010????????  :  Instruction = "vlse8.v,e64,m1";
	    34'b0000111???????101?01100010????????  :  Instruction = "vlse16.v,e64,m1";
	    34'b0000111???????110?01100010????????  :  Instruction = "vlse32.v,e64,m1";
	    34'b0000111???????111?01100010????????  :  Instruction = "vlse64.v,e64,m1";
	    34'b0000111???????000?01100110????????  :  Instruction = "vlse8.v,e64,m2";
	    34'b0000111???????101?01100110????????  :  Instruction = "vlse16.v,e64,m2";
	    34'b0000111???????110?01100110????????  :  Instruction = "vlse32.v,e64,m2";
	    34'b0000111???????111?01100110????????  :  Instruction = "vlse64.v,e64,m2";
	    34'b0000111???????000?01101010????????  :  Instruction = "vlse8.v,e64,m4";
	    34'b0000111???????101?01101010????????  :  Instruction = "vlse16.v,e64,m4";
	    34'b0000111???????110?01101010????????  :  Instruction = "vlse32.v,e64,m4";
	    34'b0000111???????111?01101010????????  :  Instruction = "vlse64.v,e64,m4";
	    34'b0000111???????000?01101110????????  :  Instruction = "vlse8.v,e64,m8";
	    34'b0000111???????101?01101110????????  :  Instruction = "vlse16.v,e64,m8";
	    34'b0000111???????110?01101110????????  :  Instruction = "vlse32.v,e64,m8";
	    34'b0000111???????111?01101110????????  :  Instruction = "vlse64.v,e64,m8";
	    34'b0000111???????111?011101?1????????  :  Instruction = "vl[uo]xei64.v,e64,mf8";
	    34'b0000111???????110?011110?1????????  :  Instruction = "vl[uo]xei32.v,e64,mf4";
	    34'b0000111???????111?011110?1????????  :  Instruction = "vl[uo]xei64.v,e64,mf4";
	    34'b0000111???????101?011111?1????????  :  Instruction = "vl[uo]xei16.v,e64,mf2";
	    34'b0000111???????110?011111?1????????  :  Instruction = "vl[uo]xei32.v,e64,mf2";
	    34'b0000111???????111?011111?1????????  :  Instruction = "vl[uo]xei64.v,e64,mf2";
	    34'b0000111???????000?011000?1????????  :  Instruction = "vl[uo]xei8.v,e64,m1";
	    34'b0000111???????101?011000?1????????  :  Instruction = "vl[uo]xei16.v,e64,m1";
	    34'b0000111???????110?011000?1????????  :  Instruction = "vl[uo]xei32.v,e64,m1";
	    34'b0000111???????111?011000?1????????  :  Instruction = "vl[uo]xei64.v,e64,m1";
	    34'b0000111???????000?011001?1????????  :  Instruction = "vl[uo]xei8.v,e64,m2";
	    34'b0000111???????101?011001?1????????  :  Instruction = "vl[uo]xei16.v,e64,m2";
	    34'b0000111???????110?011001?1????????  :  Instruction = "vl[uo]xei32.v,e64,m2";
	    34'b0000111???????111?011001?1????????  :  Instruction = "vl[uo]xei64.v,e64,m2";
	    34'b0000111???????000?011010?1????????  :  Instruction = "vl[uo]xei8.v,e64,m4";
	    34'b0000111???????101?011010?1????????  :  Instruction = "vl[uo]xei16.v,e64,m4";
	    34'b0000111???????110?011010?1????????  :  Instruction = "vl[uo]xei32.v,e64,m4";
	    34'b0000111???????111?011010?1????????  :  Instruction = "vl[uo]xei64.v,e64,m4";
	    34'b0000111???????000?011011?1????????  :  Instruction = "vl[uo]xei8.v,e64,m8";
	    34'b0000111???????101?011011?1????????  :  Instruction = "vl[uo]xei16.v,e64,m8";
	    34'b0000111???????110?011011?1????????  :  Instruction = "vl[uo]xei32.v,e64,m8";
	    34'b0000111???????111?011011?1????????  :  Instruction = "vl[uo]xei64.v,e64,m8";
	    34'b0000111???????111?01110100?0000001  :  Instruction = "vlseg2e64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000001  :  Instruction = "vlseg2e32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000001  :  Instruction = "vlseg2e64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000001  :  Instruction = "vlseg2e16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000001  :  Instruction = "vlseg2e32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000001  :  Instruction = "vlseg2e64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000001  :  Instruction = "vlseg2e8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000001  :  Instruction = "vlseg2e16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000001  :  Instruction = "vlseg2e32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000001  :  Instruction = "vlseg2e64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000001  :  Instruction = "vlseg2e8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000001  :  Instruction = "vlseg2e16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000001  :  Instruction = "vlseg2e32[ff].v,e64,m2";
	    34'b0000111???????111?01100100?0000001  :  Instruction = "vlseg2e64[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000001  :  Instruction = "vlseg2e8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000001  :  Instruction = "vlseg2e16[ff].v,e64,m4";
	    34'b0000111???????110?01101000?0000001  :  Instruction = "vlseg2e32[ff].v,e64,m4";
	    34'b0000111???????111?01101000?0000001  :  Instruction = "vlseg2e64[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000001  :  Instruction = "vlseg2e8[ff].v,e64,m8";
	    34'b0000111???????101?01101100?0000001  :  Instruction = "vlseg2e16[ff].v,e64,m8";
	    34'b0000111???????110?01101100?0000001  :  Instruction = "vlseg2e32[ff].v,e64,m8";
	    34'b0000111???????111?01101100?0000001  :  Instruction = "vlseg2e64[ff].v,e64,m8";
	    34'b0000111???????000?011???0001000001  :  Instruction = "vl2re8.v,e64";
	    34'b0000111???????101?011???0001000001  :  Instruction = "vl2re16.v,e64";
	    34'b0000111???????110?011???0001000001  :  Instruction = "vl2re32.v,e64";
	    34'b0000111???????111?011???0001000001  :  Instruction = "vl2re64.v,e64";
	    34'b0000111???????111?01110110?????001  :  Instruction = "vlsseg2e64.v,e64,mf8";
	    34'b0000111???????110?01111010?????001  :  Instruction = "vlsseg2e32.v,e64,mf4";
	    34'b0000111???????111?01111010?????001  :  Instruction = "vlsseg2e64.v,e64,mf4";
	    34'b0000111???????101?01111110?????001  :  Instruction = "vlsseg2e16.v,e64,mf2";
	    34'b0000111???????110?01111110?????001  :  Instruction = "vlsseg2e32.v,e64,mf2";
	    34'b0000111???????111?01111110?????001  :  Instruction = "vlsseg2e64.v,e64,mf2";
	    34'b0000111???????000?01100010?????001  :  Instruction = "vlsseg2e8.v,e64,m1";
	    34'b0000111???????101?01100010?????001  :  Instruction = "vlsseg2e16.v,e64,m1";
	    34'b0000111???????110?01100010?????001  :  Instruction = "vlsseg2e32.v,e64,m1";
	    34'b0000111???????111?01100010?????001  :  Instruction = "vlsseg2e64.v,e64,m1";
	    34'b0000111???????000?01100110?????001  :  Instruction = "vlsseg2e8.v,e64,m2";
	    34'b0000111???????101?01100110?????001  :  Instruction = "vlsseg2e16.v,e64,m2";
	    34'b0000111???????110?01100110?????001  :  Instruction = "vlsseg2e32.v,e64,m2";
	    34'b0000111???????111?01100110?????001  :  Instruction = "vlsseg2e64.v,e64,m2";
	    34'b0000111???????000?01101010?????001  :  Instruction = "vlsseg2e8.v,e64,m4";
	    34'b0000111???????101?01101010?????001  :  Instruction = "vlsseg2e16.v,e64,m4";
	    34'b0000111???????110?01101010?????001  :  Instruction = "vlsseg2e32.v,e64,m4";
	    34'b0000111???????111?01101010?????001  :  Instruction = "vlsseg2e64.v,e64,m4";
	    34'b0000111???????000?01101110?????001  :  Instruction = "vlsseg2e8.v,e64,m8";
	    34'b0000111???????101?01101110?????001  :  Instruction = "vlsseg2e16.v,e64,m8";
	    34'b0000111???????110?01101110?????001  :  Instruction = "vlsseg2e32.v,e64,m8";
	    34'b0000111???????111?011101?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e64,mf8";
	    34'b0000111???????110?011110?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e64,mf4";
	    34'b0000111???????111?011110?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e64,mf4";
	    34'b0000111???????101?011111?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e64,mf2";
	    34'b0000111???????110?011111?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e64,mf2";
	    34'b0000111???????111?011111?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e64,mf2";
	    34'b0000111???????000?011000?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e64,m1";
	    34'b0000111???????101?011000?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e64,m1";
	    34'b0000111???????110?011000?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e64,m1";
	    34'b0000111???????111?011000?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e64,m1";
	    34'b0000111???????000?011001?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e64,m2";
	    34'b0000111???????101?011001?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e64,m2";
	    34'b0000111???????110?011001?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e64,m2";
	    34'b0000111???????111?011001?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e64,m2";
	    34'b0000111???????000?011010?1?????001  :  Instruction = "vl[uo]xseg2ei8.v,e64,m4";
	    34'b0000111???????101?011010?1?????001  :  Instruction = "vl[uo]xseg2ei16.v,e64,m4";
	    34'b0000111???????110?011010?1?????001  :  Instruction = "vl[uo]xseg2ei32.v,e64,m4";
	    34'b0000111???????111?011010?1?????001  :  Instruction = "vl[uo]xseg2ei64.v,e64,m4";
	    34'b0000111???????111?01110100?0000010  :  Instruction = "vlseg3e64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000010  :  Instruction = "vlseg3e32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000010  :  Instruction = "vlseg3e64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000010  :  Instruction = "vlseg3e16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000010  :  Instruction = "vlseg3e32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000010  :  Instruction = "vlseg3e64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000010  :  Instruction = "vlseg3e8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000010  :  Instruction = "vlseg3e16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000010  :  Instruction = "vlseg3e32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000010  :  Instruction = "vlseg3e64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000010  :  Instruction = "vlseg3e8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000010  :  Instruction = "vlseg3e16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000010  :  Instruction = "vlseg3e32[ff].v,e64,m2";
	    34'b0000111???????111?01100100?0000010  :  Instruction = "vlseg3e64[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000010  :  Instruction = "vlseg3e8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000010  :  Instruction = "vlseg3e16[ff].v,e64,m4";
	    34'b0000111???????110?01101000?0000010  :  Instruction = "vlseg3e32[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000010  :  Instruction = "vlseg3e8[ff].v,e64,m8";
	    34'b0000111???????101?01101100?0000010  :  Instruction = "vlseg3e16[ff].v,e64,m8";
	    34'b0000111???????111?01110110?????010  :  Instruction = "vlsseg3e64.v,e64,mf8";
	    34'b0000111???????110?01111010?????010  :  Instruction = "vlsseg3e32.v,e64,mf4";
	    34'b0000111???????111?01111010?????010  :  Instruction = "vlsseg3e64.v,e64,mf4";
	    34'b0000111???????101?01111110?????010  :  Instruction = "vlsseg3e16.v,e64,mf2";
	    34'b0000111???????110?01111110?????010  :  Instruction = "vlsseg3e32.v,e64,mf2";
	    34'b0000111???????111?01111110?????010  :  Instruction = "vlsseg3e64.v,e64,mf2";
	    34'b0000111???????000?01100010?????010  :  Instruction = "vlsseg3e8.v,e64,m1";
	    34'b0000111???????101?01100010?????010  :  Instruction = "vlsseg3e16.v,e64,m1";
	    34'b0000111???????110?01100010?????010  :  Instruction = "vlsseg3e32.v,e64,m1";
	    34'b0000111???????111?01100010?????010  :  Instruction = "vlsseg3e64.v,e64,m1";
	    34'b0000111???????000?01100110?????010  :  Instruction = "vlsseg3e8.v,e64,m2";
	    34'b0000111???????101?01100110?????010  :  Instruction = "vlsseg3e16.v,e64,m2";
	    34'b0000111???????110?01100110?????010  :  Instruction = "vlsseg3e32.v,e64,m2";
	    34'b0000111???????111?01100110?????010  :  Instruction = "vlsseg3e64.v,e64,m2";
	    34'b0000111???????000?01101010?????010  :  Instruction = "vlsseg3e8.v,e64,m4";
	    34'b0000111???????101?01101010?????010  :  Instruction = "vlsseg3e16.v,e64,m4";
	    34'b0000111???????110?01101010?????010  :  Instruction = "vlsseg3e32.v,e64,m4";
	    34'b0000111???????000?01101110?????010  :  Instruction = "vlsseg3e8.v,e64,m8";
	    34'b0000111???????101?01101110?????010  :  Instruction = "vlsseg3e16.v,e64,m8";
	    34'b0000111???????111?011101?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e64,mf8";
	    34'b0000111???????110?011110?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e64,mf4";
	    34'b0000111???????111?011110?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e64,mf4";
	    34'b0000111???????101?011111?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e64,mf2";
	    34'b0000111???????110?011111?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e64,mf2";
	    34'b0000111???????111?011111?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e64,mf2";
	    34'b0000111???????000?011000?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e64,m1";
	    34'b0000111???????101?011000?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e64,m1";
	    34'b0000111???????110?011000?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e64,m1";
	    34'b0000111???????111?011000?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e64,m1";
	    34'b0000111???????000?011001?1?????010  :  Instruction = "vl[uo]xseg3ei8.v,e64,m2";
	    34'b0000111???????101?011001?1?????010  :  Instruction = "vl[uo]xseg3ei16.v,e64,m2";
	    34'b0000111???????110?011001?1?????010  :  Instruction = "vl[uo]xseg3ei32.v,e64,m2";
	    34'b0000111???????111?011001?1?????010  :  Instruction = "vl[uo]xseg3ei64.v,e64,m2";
	    34'b0000111???????111?01110100?0000011  :  Instruction = "vlseg4e64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000011  :  Instruction = "vlseg4e32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000011  :  Instruction = "vlseg4e64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000011  :  Instruction = "vlseg4e16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000011  :  Instruction = "vlseg4e32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000011  :  Instruction = "vlseg4e64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000011  :  Instruction = "vlseg4e8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000011  :  Instruction = "vlseg4e16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000011  :  Instruction = "vlseg4e32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000011  :  Instruction = "vlseg4e64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000011  :  Instruction = "vlseg4e8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000011  :  Instruction = "vlseg4e16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000011  :  Instruction = "vlseg4e32[ff].v,e64,m2";
	    34'b0000111???????111?01100100?0000011  :  Instruction = "vlseg4e64[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000011  :  Instruction = "vlseg4e8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000011  :  Instruction = "vlseg4e16[ff].v,e64,m4";
	    34'b0000111???????110?01101000?0000011  :  Instruction = "vlseg4e32[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000011  :  Instruction = "vlseg4e8[ff].v,e64,m8";
	    34'b0000111???????101?01101100?0000011  :  Instruction = "vlseg4e16[ff].v,e64,m8";
	    34'b0000111???????111?01110110?????011  :  Instruction = "vlsseg4e64.v,e64,mf8";
	    34'b0000111???????110?01111010?????011  :  Instruction = "vlsseg4e32.v,e64,mf4";
	    34'b0000111???????111?01111010?????011  :  Instruction = "vlsseg4e64.v,e64,mf4";
	    34'b0000111???????101?01111110?????011  :  Instruction = "vlsseg4e16.v,e64,mf2";
	    34'b0000111???????110?01111110?????011  :  Instruction = "vlsseg4e32.v,e64,mf2";
	    34'b0000111???????111?01111110?????011  :  Instruction = "vlsseg4e64.v,e64,mf2";
	    34'b0000111???????000?01100010?????011  :  Instruction = "vlsseg4e8.v,e64,m1";
	    34'b0000111???????101?01100010?????011  :  Instruction = "vlsseg4e16.v,e64,m1";
	    34'b0000111???????110?01100010?????011  :  Instruction = "vlsseg4e32.v,e64,m1";
	    34'b0000111???????111?01100010?????011  :  Instruction = "vlsseg4e64.v,e64,m1";
	    34'b0000111???????000?01100110?????011  :  Instruction = "vlsseg4e8.v,e64,m2";
	    34'b0000111???????101?01100110?????011  :  Instruction = "vlsseg4e16.v,e64,m2";
	    34'b0000111???????110?01100110?????011  :  Instruction = "vlsseg4e32.v,e64,m2";
	    34'b0000111???????111?01100110?????011  :  Instruction = "vlsseg4e64.v,e64,m2";
	    34'b0000111???????000?01101010?????011  :  Instruction = "vlsseg4e8.v,e64,m4";
	    34'b0000111???????101?01101010?????011  :  Instruction = "vlsseg4e16.v,e64,m4";
	    34'b0000111???????110?01101010?????011  :  Instruction = "vlsseg4e32.v,e64,m4";
	    34'b0000111???????000?01101110?????011  :  Instruction = "vlsseg4e8.v,e64,m8";
	    34'b0000111???????101?01101110?????011  :  Instruction = "vlsseg4e16.v,e64,m8";
	    34'b0000111???????000?011???0001000011  :  Instruction = "vl4re8.v,e64";
	    34'b0000111???????101?011???0001000011  :  Instruction = "vl4re16.v,e64";
	    34'b0000111???????110?011???0001000011  :  Instruction = "vl4re32.v,e64";
	    34'b0000111???????111?011???0001000011  :  Instruction = "vl4re64.v,e64";
	    34'b0000111???????111?011101?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e64,mf8";
	    34'b0000111???????110?011110?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e64,mf4";
	    34'b0000111???????111?011110?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e64,mf4";
	    34'b0000111???????101?011111?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e64,mf2";
	    34'b0000111???????110?011111?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e64,mf2";
	    34'b0000111???????111?011111?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e64,mf2";
	    34'b0000111???????000?011000?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e64,m1";
	    34'b0000111???????101?011000?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e64,m1";
	    34'b0000111???????110?011000?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e64,m1";
	    34'b0000111???????111?011000?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e64,m1";
	    34'b0000111???????000?011001?1?????011  :  Instruction = "vl[uo]xseg4ei8.v,e64,m2";
	    34'b0000111???????101?011001?1?????011  :  Instruction = "vl[uo]xseg4ei16.v,e64,m2";
	    34'b0000111???????110?011001?1?????011  :  Instruction = "vl[uo]xseg4ei32.v,e64,m2";
	    34'b0000111???????111?011001?1?????011  :  Instruction = "vl[uo]xseg4ei64.v,e64,m2";
	    34'b0000111???????111?01110100?0000100  :  Instruction = "vlseg5e64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000100  :  Instruction = "vlseg5e32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000100  :  Instruction = "vlseg5e64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000100  :  Instruction = "vlseg5e16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000100  :  Instruction = "vlseg5e32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000100  :  Instruction = "vlseg5e64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000100  :  Instruction = "vlseg5e8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000100  :  Instruction = "vlseg5e16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000100  :  Instruction = "vlseg5e32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000100  :  Instruction = "vlseg5e64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000100  :  Instruction = "vlseg5e8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000100  :  Instruction = "vlseg5e16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000100  :  Instruction = "vlseg5e32[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000100  :  Instruction = "vlseg5e8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000100  :  Instruction = "vlseg5e16[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000100  :  Instruction = "vlseg5e8[ff].v,e64,m8";
	    34'b0000111???????111?01110110?????100  :  Instruction = "vlsseg5e64.v,e64,mf8";
	    34'b0000111???????110?01111010?????100  :  Instruction = "vlsseg5e32.v,e64,mf4";
	    34'b0000111???????111?01111010?????100  :  Instruction = "vlsseg5e64.v,e64,mf4";
	    34'b0000111???????101?01111110?????100  :  Instruction = "vlsseg5e16.v,e64,mf2";
	    34'b0000111???????110?01111110?????100  :  Instruction = "vlsseg5e32.v,e64,mf2";
	    34'b0000111???????111?01111110?????100  :  Instruction = "vlsseg5e64.v,e64,mf2";
	    34'b0000111???????000?01100010?????100  :  Instruction = "vlsseg5e8.v,e64,m1";
	    34'b0000111???????101?01100010?????100  :  Instruction = "vlsseg5e16.v,e64,m1";
	    34'b0000111???????110?01100010?????100  :  Instruction = "vlsseg5e32.v,e64,m1";
	    34'b0000111???????111?01100010?????100  :  Instruction = "vlsseg5e64.v,e64,m1";
	    34'b0000111???????000?01100110?????100  :  Instruction = "vlsseg5e8.v,e64,m2";
	    34'b0000111???????101?01100110?????100  :  Instruction = "vlsseg5e16.v,e64,m2";
	    34'b0000111???????110?01100110?????100  :  Instruction = "vlsseg5e32.v,e64,m2";
	    34'b0000111???????000?01101010?????100  :  Instruction = "vlsseg5e8.v,e64,m4";
	    34'b0000111???????101?01101010?????100  :  Instruction = "vlsseg5e16.v,e64,m4";
	    34'b0000111???????000?01101110?????100  :  Instruction = "vlsseg5e8.v,e64,m8";
	    34'b0000111???????111?011101?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e64,mf8";
	    34'b0000111???????110?011110?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e64,mf4";
	    34'b0000111???????111?011110?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e64,mf4";
	    34'b0000111???????101?011111?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e64,mf2";
	    34'b0000111???????110?011111?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e64,mf2";
	    34'b0000111???????111?011111?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e64,mf2";
	    34'b0000111???????000?011000?1?????100  :  Instruction = "vl[uo]xseg5ei8.v,e64,m1";
	    34'b0000111???????101?011000?1?????100  :  Instruction = "vl[uo]xseg5ei16.v,e64,m1";
	    34'b0000111???????110?011000?1?????100  :  Instruction = "vl[uo]xseg5ei32.v,e64,m1";
	    34'b0000111???????111?011000?1?????100  :  Instruction = "vl[uo]xseg5ei64.v,e64,m1";
	    34'b0000111???????111?01110100?0000101  :  Instruction = "vlseg6e64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000101  :  Instruction = "vlseg6e32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000101  :  Instruction = "vlseg6e64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000101  :  Instruction = "vlseg6e16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000101  :  Instruction = "vlseg6e32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000101  :  Instruction = "vlseg6e64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000101  :  Instruction = "vlseg6e8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000101  :  Instruction = "vlseg6e16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000101  :  Instruction = "vlseg6e32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000101  :  Instruction = "vlseg6e64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000101  :  Instruction = "vlseg6e8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000101  :  Instruction = "vlseg6e16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000101  :  Instruction = "vlseg6e32[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000101  :  Instruction = "vlseg6e8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000101  :  Instruction = "vlseg6e16[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000101  :  Instruction = "vlseg6e8[ff].v,e64,m8";
	    34'b0000111???????111?01110110?????101  :  Instruction = "vlsseg6e64.v,e64,mf8";
	    34'b0000111???????110?01111010?????101  :  Instruction = "vlsseg6e32.v,e64,mf4";
	    34'b0000111???????111?01111010?????101  :  Instruction = "vlsseg6e64.v,e64,mf4";
	    34'b0000111???????101?01111110?????101  :  Instruction = "vlsseg6e16.v,e64,mf2";
	    34'b0000111???????110?01111110?????101  :  Instruction = "vlsseg6e32.v,e64,mf2";
	    34'b0000111???????111?01111110?????101  :  Instruction = "vlsseg6e64.v,e64,mf2";
	    34'b0000111???????000?01100010?????101  :  Instruction = "vlsseg6e8.v,e64,m1";
	    34'b0000111???????101?01100010?????101  :  Instruction = "vlsseg6e16.v,e64,m1";
	    34'b0000111???????110?01100010?????101  :  Instruction = "vlsseg6e32.v,e64,m1";
	    34'b0000111???????111?01100010?????101  :  Instruction = "vlsseg6e64.v,e64,m1";
	    34'b0000111???????000?01100110?????101  :  Instruction = "vlsseg6e8.v,e64,m2";
	    34'b0000111???????101?01100110?????101  :  Instruction = "vlsseg6e16.v,e64,m2";
	    34'b0000111???????110?01100110?????101  :  Instruction = "vlsseg6e32.v,e64,m2";
	    34'b0000111???????000?01101010?????101  :  Instruction = "vlsseg6e8.v,e64,m4";
	    34'b0000111???????101?01101010?????101  :  Instruction = "vlsseg6e16.v,e64,m4";
	    34'b0000111???????000?01101110?????101  :  Instruction = "vlsseg6e8.v,e64,m8";
	    34'b0000111???????111?011101?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e64,mf8";
	    34'b0000111???????110?011110?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e64,mf4";
	    34'b0000111???????111?011110?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e64,mf4";
	    34'b0000111???????101?011111?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e64,mf2";
	    34'b0000111???????110?011111?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e64,mf2";
	    34'b0000111???????111?011111?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e64,mf2";
	    34'b0000111???????000?011000?1?????101  :  Instruction = "vl[uo]xseg6ei8.v,e64,m1";
	    34'b0000111???????101?011000?1?????101  :  Instruction = "vl[uo]xseg6ei16.v,e64,m1";
	    34'b0000111???????110?011000?1?????101  :  Instruction = "vl[uo]xseg6ei32.v,e64,m1";
	    34'b0000111???????111?011000?1?????101  :  Instruction = "vl[uo]xseg6ei64.v,e64,m1";
	    34'b0000111???????111?01110100?0000110  :  Instruction = "vlseg7e64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000110  :  Instruction = "vlseg7e32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000110  :  Instruction = "vlseg7e64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000110  :  Instruction = "vlseg7e16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000110  :  Instruction = "vlseg7e32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000110  :  Instruction = "vlseg7e64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000110  :  Instruction = "vlseg7e8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000110  :  Instruction = "vlseg7e16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000110  :  Instruction = "vlseg7e32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000110  :  Instruction = "vlseg7e64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000110  :  Instruction = "vlseg7e8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000110  :  Instruction = "vlseg7e16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000110  :  Instruction = "vlseg7e32[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000110  :  Instruction = "vlseg7e8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000110  :  Instruction = "vlseg7e16[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000110  :  Instruction = "vlseg7e8[ff].v,e64,m8";
	    34'b0000111???????111?01110110?????110  :  Instruction = "vlsseg7e64.v,e64,mf8";
	    34'b0000111???????110?01111010?????110  :  Instruction = "vlsseg7e32.v,e64,mf4";
	    34'b0000111???????111?01111010?????110  :  Instruction = "vlsseg7e64.v,e64,mf4";
	    34'b0000111???????101?01111110?????110  :  Instruction = "vlsseg7e16.v,e64,mf2";
	    34'b0000111???????110?01111110?????110  :  Instruction = "vlsseg7e32.v,e64,mf2";
	    34'b0000111???????111?01111110?????110  :  Instruction = "vlsseg7e64.v,e64,mf2";
	    34'b0000111???????000?01100010?????110  :  Instruction = "vlsseg7e8.v,e64,m1";
	    34'b0000111???????101?01100010?????110  :  Instruction = "vlsseg7e16.v,e64,m1";
	    34'b0000111???????110?01100010?????110  :  Instruction = "vlsseg7e32.v,e64,m1";
	    34'b0000111???????111?01100010?????110  :  Instruction = "vlsseg7e64.v,e64,m1";
	    34'b0000111???????000?01100110?????110  :  Instruction = "vlsseg7e8.v,e64,m2";
	    34'b0000111???????101?01100110?????110  :  Instruction = "vlsseg7e16.v,e64,m2";
	    34'b0000111???????110?01100110?????110  :  Instruction = "vlsseg7e32.v,e64,m2";
	    34'b0000111???????000?01101010?????110  :  Instruction = "vlsseg7e8.v,e64,m4";
	    34'b0000111???????101?01101010?????110  :  Instruction = "vlsseg7e16.v,e64,m4";
	    34'b0000111???????000?01101110?????110  :  Instruction = "vlsseg7e8.v,e64,m8";
	    34'b0000111???????111?011101?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e64,mf8";
	    34'b0000111???????110?011110?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e64,mf4";
	    34'b0000111???????111?011110?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e64,mf4";
	    34'b0000111???????101?011111?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e64,mf2";
	    34'b0000111???????110?011111?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e64,mf2";
	    34'b0000111???????111?011111?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e64,mf2";
	    34'b0000111???????000?011000?1?????110  :  Instruction = "vl[uo]xseg7ei8.v,e64,m1";
	    34'b0000111???????101?011000?1?????110  :  Instruction = "vl[uo]xseg7ei16.v,e64,m1";
	    34'b0000111???????110?011000?1?????110  :  Instruction = "vl[uo]xseg7ei32.v,e64,m1";
	    34'b0000111???????111?011000?1?????110  :  Instruction = "vl[uo]xseg7ei64.v,e64,m1";
	    34'b0000111???????111?01110100?0000111  :  Instruction = "vlseg8e64[ff].v,e64,mf8";
	    34'b0000111???????110?01111000?0000111  :  Instruction = "vlseg8e32[ff].v,e64,mf4";
	    34'b0000111???????111?01111000?0000111  :  Instruction = "vlseg8e64[ff].v,e64,mf4";
	    34'b0000111???????101?01111100?0000111  :  Instruction = "vlseg8e16[ff].v,e64,mf2";
	    34'b0000111???????110?01111100?0000111  :  Instruction = "vlseg8e32[ff].v,e64,mf2";
	    34'b0000111???????111?01111100?0000111  :  Instruction = "vlseg8e64[ff].v,e64,mf2";
	    34'b0000111???????000?01100000?0000111  :  Instruction = "vlseg8e8[ff].v,e64,m1";
	    34'b0000111???????101?01100000?0000111  :  Instruction = "vlseg8e16[ff].v,e64,m1";
	    34'b0000111???????110?01100000?0000111  :  Instruction = "vlseg8e32[ff].v,e64,m1";
	    34'b0000111???????111?01100000?0000111  :  Instruction = "vlseg8e64[ff].v,e64,m1";
	    34'b0000111???????000?01100100?0000111  :  Instruction = "vlseg8e8[ff].v,e64,m2";
	    34'b0000111???????101?01100100?0000111  :  Instruction = "vlseg8e16[ff].v,e64,m2";
	    34'b0000111???????110?01100100?0000111  :  Instruction = "vlseg8e32[ff].v,e64,m2";
	    34'b0000111???????000?01101000?0000111  :  Instruction = "vlseg8e8[ff].v,e64,m4";
	    34'b0000111???????101?01101000?0000111  :  Instruction = "vlseg8e16[ff].v,e64,m4";
	    34'b0000111???????000?01101100?0000111  :  Instruction = "vlseg8e8[ff].v,e64,m8";
	    34'b0000111???????000?011???0001000111  :  Instruction = "vl8re8.v,e64";
	    34'b0000111???????101?011???0001000111  :  Instruction = "vl8re16.v,e64";
	    34'b0000111???????110?011???0001000111  :  Instruction = "vl8re32.v,e64";
	    34'b0000111???????111?011???0001000111  :  Instruction = "vl8re64.v,e64";
	    34'b0000111???????111?01110110?????111  :  Instruction = "vlsseg8e64.v,e64,mf8";
	    34'b0000111???????110?01111010?????111  :  Instruction = "vlsseg8e32.v,e64,mf4";
	    34'b0000111???????111?01111010?????111  :  Instruction = "vlsseg8e64.v,e64,mf4";
	    34'b0000111???????101?01111110?????111  :  Instruction = "vlsseg8e16.v,e64,mf2";
	    34'b0000111???????110?01111110?????111  :  Instruction = "vlsseg8e32.v,e64,mf2";
	    34'b0000111???????111?01111110?????111  :  Instruction = "vlsseg8e64.v,e64,mf2";
	    34'b0000111???????000?01100010?????111  :  Instruction = "vlsseg8e8.v,e64,m1";
	    34'b0000111???????101?01100010?????111  :  Instruction = "vlsseg8e16.v,e64,m1";
	    34'b0000111???????110?01100010?????111  :  Instruction = "vlsseg8e32.v,e64,m1";
	    34'b0000111???????111?01100010?????111  :  Instruction = "vlsseg8e64.v,e64,m1";
	    34'b0000111???????000?01100110?????111  :  Instruction = "vlsseg8e8.v,e64,m2";
	    34'b0000111???????101?01100110?????111  :  Instruction = "vlsseg8e16.v,e64,m2";
	    34'b0000111???????110?01100110?????111  :  Instruction = "vlsseg8e32.v,e64,m2";
	    34'b0000111???????000?01101010?????111  :  Instruction = "vlsseg8e8.v,e64,m4";
	    34'b0000111???????101?01101010?????111  :  Instruction = "vlsseg8e16.v,e64,m4";
	    34'b0000111???????000?01101110?????111  :  Instruction = "vlsseg8e8.v,e64,m8";
	    34'b0000111???????111?011101?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e64,mf8";
	    34'b0000111???????110?011110?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e64,mf4";
	    34'b0000111???????111?011110?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e64,mf4";
	    34'b0000111???????101?011111?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e64,mf2";
	    34'b0000111???????110?011111?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e64,mf2";
	    34'b0000111???????111?011111?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e64,mf2";
	    34'b0000111???????000?011000?1?????111  :  Instruction = "vl[uo]xseg8ei8.v,e64,m1";
	    34'b0000111???????101?011000?1?????111  :  Instruction = "vl[uo]xseg8ei16.v,e64,m1";
	    34'b0000111???????110?011000?1?????111  :  Instruction = "vl[uo]xseg8ei32.v,e64,m1";
	    34'b0000111???????111?011000?1?????111  :  Instruction = "vl[uo]xseg8ei64.v,e64,m1";
	    34'b0100111???????111?01110100?0000???  :  Instruction = "vse64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000???  :  Instruction = "vse32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000???  :  Instruction = "vse64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000???  :  Instruction = "vse16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000???  :  Instruction = "vse32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000???  :  Instruction = "vse64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000???  :  Instruction = "vse8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000???  :  Instruction = "vse16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000???  :  Instruction = "vse32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000???  :  Instruction = "vse64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000???  :  Instruction = "vse8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000???  :  Instruction = "vse16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000???  :  Instruction = "vse32[ff].v,e64,m2";
	    34'b0100111???????111?01100100?0000???  :  Instruction = "vse64[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000???  :  Instruction = "vse8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000???  :  Instruction = "vse16[ff].v,e64,m4";
	    34'b0100111???????110?01101000?0000???  :  Instruction = "vse32[ff].v,e64,m4";
	    34'b0100111???????111?01101000?0000???  :  Instruction = "vse64[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000???  :  Instruction = "vse8[ff].v,e64,m8";
	    34'b0100111???????101?01101100?0000???  :  Instruction = "vse16[ff].v,e64,m8";
	    34'b0100111???????110?01101100?0000???  :  Instruction = "vse32[ff].v,e64,m8";
	    34'b0100111???????111?01101100?0000???  :  Instruction = "vse64[ff].v,e64,m8";
	    34'b0100111???????000?011???0001000000  :  Instruction = "vs1r.v,e64";
	    34'b0100111???????111?01110110????????  :  Instruction = "vsse64.v,e64,mf8";
	    34'b0100111???????110?01111010????????  :  Instruction = "vsse32.v,e64,mf4";
	    34'b0100111???????111?01111010????????  :  Instruction = "vsse64.v,e64,mf4";
	    34'b0100111???????101?01111110????????  :  Instruction = "vsse16.v,e64,mf2";
	    34'b0100111???????110?01111110????????  :  Instruction = "vsse32.v,e64,mf2";
	    34'b0100111???????111?01111110????????  :  Instruction = "vsse64.v,e64,mf2";
	    34'b0100111???????000?01100010????????  :  Instruction = "vsse8.v,e64,m1";
	    34'b0100111???????101?01100010????????  :  Instruction = "vsse16.v,e64,m1";
	    34'b0100111???????110?01100010????????  :  Instruction = "vsse32.v,e64,m1";
	    34'b0100111???????111?01100010????????  :  Instruction = "vsse64.v,e64,m1";
	    34'b0100111???????000?01100110????????  :  Instruction = "vsse8.v,e64,m2";
	    34'b0100111???????101?01100110????????  :  Instruction = "vsse16.v,e64,m2";
	    34'b0100111???????110?01100110????????  :  Instruction = "vsse32.v,e64,m2";
	    34'b0100111???????111?01100110????????  :  Instruction = "vsse64.v,e64,m2";
	    34'b0100111???????000?01101010????????  :  Instruction = "vsse8.v,e64,m4";
	    34'b0100111???????101?01101010????????  :  Instruction = "vsse16.v,e64,m4";
	    34'b0100111???????110?01101010????????  :  Instruction = "vsse32.v,e64,m4";
	    34'b0100111???????111?01101010????????  :  Instruction = "vsse64.v,e64,m4";
	    34'b0100111???????000?01101110????????  :  Instruction = "vsse8.v,e64,m8";
	    34'b0100111???????101?01101110????????  :  Instruction = "vsse16.v,e64,m8";
	    34'b0100111???????110?01101110????????  :  Instruction = "vsse32.v,e64,m8";
	    34'b0100111???????111?01101110????????  :  Instruction = "vsse64.v,e64,m8";
	    34'b0100111???????111?011101?1????????  :  Instruction = "vs[uo]xei64.v,e64,mf8";
	    34'b0100111???????110?011110?1????????  :  Instruction = "vs[uo]xei32.v,e64,mf4";
	    34'b0100111???????111?011110?1????????  :  Instruction = "vs[uo]xei64.v,e64,mf4";
	    34'b0100111???????101?011111?1????????  :  Instruction = "vs[uo]xei16.v,e64,mf2";
	    34'b0100111???????110?011111?1????????  :  Instruction = "vs[uo]xei32.v,e64,mf2";
	    34'b0100111???????111?011111?1????????  :  Instruction = "vs[uo]xei64.v,e64,mf2";
	    34'b0100111???????000?011000?1????????  :  Instruction = "vs[uo]xei8.v,e64,m1";
	    34'b0100111???????101?011000?1????????  :  Instruction = "vs[uo]xei16.v,e64,m1";
	    34'b0100111???????110?011000?1????????  :  Instruction = "vs[uo]xei32.v,e64,m1";
	    34'b0100111???????111?011000?1????????  :  Instruction = "vs[uo]xei64.v,e64,m1";
	    34'b0100111???????000?011001?1????????  :  Instruction = "vs[uo]xei8.v,e64,m2";
	    34'b0100111???????101?011001?1????????  :  Instruction = "vs[uo]xei16.v,e64,m2";
	    34'b0100111???????110?011001?1????????  :  Instruction = "vs[uo]xei32.v,e64,m2";
	    34'b0100111???????111?011001?1????????  :  Instruction = "vs[uo]xei64.v,e64,m2";
	    34'b0100111???????000?011010?1????????  :  Instruction = "vs[uo]xei8.v,e64,m4";
	    34'b0100111???????101?011010?1????????  :  Instruction = "vs[uo]xei16.v,e64,m4";
	    34'b0100111???????110?011010?1????????  :  Instruction = "vs[uo]xei32.v,e64,m4";
	    34'b0100111???????111?011010?1????????  :  Instruction = "vs[uo]xei64.v,e64,m4";
	    34'b0100111???????000?011011?1????????  :  Instruction = "vs[uo]xei8.v,e64,m8";
	    34'b0100111???????101?011011?1????????  :  Instruction = "vs[uo]xei16.v,e64,m8";
	    34'b0100111???????110?011011?1????????  :  Instruction = "vs[uo]xei32.v,e64,m8";
	    34'b0100111???????111?011011?1????????  :  Instruction = "vs[uo]xei64.v,e64,m8";
	    34'b0100111???????111?01110100?0000001  :  Instruction = "vsseg2e64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000001  :  Instruction = "vsseg2e32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000001  :  Instruction = "vsseg2e64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000001  :  Instruction = "vsseg2e16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000001  :  Instruction = "vsseg2e32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000001  :  Instruction = "vsseg2e64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000001  :  Instruction = "vsseg2e8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000001  :  Instruction = "vsseg2e16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000001  :  Instruction = "vsseg2e32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000001  :  Instruction = "vsseg2e64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000001  :  Instruction = "vsseg2e8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000001  :  Instruction = "vsseg2e16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000001  :  Instruction = "vsseg2e32[ff].v,e64,m2";
	    34'b0100111???????111?01100100?0000001  :  Instruction = "vsseg2e64[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000001  :  Instruction = "vsseg2e8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000001  :  Instruction = "vsseg2e16[ff].v,e64,m4";
	    34'b0100111???????110?01101000?0000001  :  Instruction = "vsseg2e32[ff].v,e64,m4";
	    34'b0100111???????111?01101000?0000001  :  Instruction = "vsseg2e64[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000001  :  Instruction = "vsseg2e8[ff].v,e64,m8";
	    34'b0100111???????101?01101100?0000001  :  Instruction = "vsseg2e16[ff].v,e64,m8";
	    34'b0100111???????110?01101100?0000001  :  Instruction = "vsseg2e32[ff].v,e64,m8";
	    34'b0100111???????000?011???0001000001  :  Instruction = "vs2r.v,e64";
	    34'b0100111???????111?01110110?????001  :  Instruction = "vssseg2e64.v,e64,mf8";
	    34'b0100111???????110?01111010?????001  :  Instruction = "vssseg2e32.v,e64,mf4";
	    34'b0100111???????111?01111010?????001  :  Instruction = "vssseg2e64.v,e64,mf4";
	    34'b0100111???????101?01111110?????001  :  Instruction = "vssseg2e16.v,e64,mf2";
	    34'b0100111???????110?01111110?????001  :  Instruction = "vssseg2e32.v,e64,mf2";
	    34'b0100111???????111?01111110?????001  :  Instruction = "vssseg2e64.v,e64,mf2";
	    34'b0100111???????000?01100010?????001  :  Instruction = "vssseg2e8.v,e64,m1";
	    34'b0100111???????101?01100010?????001  :  Instruction = "vssseg2e16.v,e64,m1";
	    34'b0100111???????110?01100010?????001  :  Instruction = "vssseg2e32.v,e64,m1";
	    34'b0100111???????111?01100010?????001  :  Instruction = "vssseg2e64.v,e64,m1";
	    34'b0100111???????000?01100110?????001  :  Instruction = "vssseg2e8.v,e64,m2";
	    34'b0100111???????101?01100110?????001  :  Instruction = "vssseg2e16.v,e64,m2";
	    34'b0100111???????110?01100110?????001  :  Instruction = "vssseg2e32.v,e64,m2";
	    34'b0100111???????111?01100110?????001  :  Instruction = "vssseg2e64.v,e64,m2";
	    34'b0100111???????000?01101010?????001  :  Instruction = "vssseg2e8.v,e64,m4";
	    34'b0100111???????101?01101010?????001  :  Instruction = "vssseg2e16.v,e64,m4";
	    34'b0100111???????110?01101010?????001  :  Instruction = "vssseg2e32.v,e64,m4";
	    34'b0100111???????111?01101010?????001  :  Instruction = "vssseg2e64.v,e64,m4";
	    34'b0100111???????000?01101110?????001  :  Instruction = "vssseg2e8.v,e64,m8";
	    34'b0100111???????101?01101110?????001  :  Instruction = "vssseg2e16.v,e64,m8";
	    34'b0100111???????110?01101110?????001  :  Instruction = "vssseg2e32.v,e64,m8";
	    34'b0100111???????111?011101?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e64,mf8";
	    34'b0100111???????110?011110?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e64,mf4";
	    34'b0100111???????111?011110?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e64,mf4";
	    34'b0100111???????101?011111?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e64,mf2";
	    34'b0100111???????110?011111?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e64,mf2";
	    34'b0100111???????111?011111?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e64,mf2";
	    34'b0100111???????000?011000?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e64,m1";
	    34'b0100111???????101?011000?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e64,m1";
	    34'b0100111???????110?011000?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e64,m1";
	    34'b0100111???????111?011000?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e64,m1";
	    34'b0100111???????000?011001?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e64,m2";
	    34'b0100111???????101?011001?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e64,m2";
	    34'b0100111???????110?011001?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e64,m2";
	    34'b0100111???????111?011001?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e64,m2";
	    34'b0100111???????000?011010?1?????001  :  Instruction = "vs[uo]xseg2ei8.v,e64,m4";
	    34'b0100111???????101?011010?1?????001  :  Instruction = "vs[uo]xseg2ei16.v,e64,m4";
	    34'b0100111???????110?011010?1?????001  :  Instruction = "vs[uo]xseg2ei32.v,e64,m4";
	    34'b0100111???????111?011010?1?????001  :  Instruction = "vs[uo]xseg2ei64.v,e64,m4";
	    34'b0100111???????111?01110100?0000010  :  Instruction = "vsseg3e64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000010  :  Instruction = "vsseg3e32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000010  :  Instruction = "vsseg3e64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000010  :  Instruction = "vsseg3e16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000010  :  Instruction = "vsseg3e32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000010  :  Instruction = "vsseg3e64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000010  :  Instruction = "vsseg3e8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000010  :  Instruction = "vsseg3e16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000010  :  Instruction = "vsseg3e32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000010  :  Instruction = "vsseg3e64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000010  :  Instruction = "vsseg3e8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000010  :  Instruction = "vsseg3e16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000010  :  Instruction = "vsseg3e32[ff].v,e64,m2";
	    34'b0100111???????111?01100100?0000010  :  Instruction = "vsseg3e64[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000010  :  Instruction = "vsseg3e8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000010  :  Instruction = "vsseg3e16[ff].v,e64,m4";
	    34'b0100111???????110?01101000?0000010  :  Instruction = "vsseg3e32[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000010  :  Instruction = "vsseg3e8[ff].v,e64,m8";
	    34'b0100111???????101?01101100?0000010  :  Instruction = "vsseg3e16[ff].v,e64,m8";
	    34'b0100111???????111?01110110?????010  :  Instruction = "vssseg3e64.v,e64,mf8";
	    34'b0100111???????110?01111010?????010  :  Instruction = "vssseg3e32.v,e64,mf4";
	    34'b0100111???????111?01111010?????010  :  Instruction = "vssseg3e64.v,e64,mf4";
	    34'b0100111???????101?01111110?????010  :  Instruction = "vssseg3e16.v,e64,mf2";
	    34'b0100111???????110?01111110?????010  :  Instruction = "vssseg3e32.v,e64,mf2";
	    34'b0100111???????111?01111110?????010  :  Instruction = "vssseg3e64.v,e64,mf2";
	    34'b0100111???????000?01100010?????010  :  Instruction = "vssseg3e8.v,e64,m1";
	    34'b0100111???????101?01100010?????010  :  Instruction = "vssseg3e16.v,e64,m1";
	    34'b0100111???????110?01100010?????010  :  Instruction = "vssseg3e32.v,e64,m1";
	    34'b0100111???????111?01100010?????010  :  Instruction = "vssseg3e64.v,e64,m1";
	    34'b0100111???????000?01100110?????010  :  Instruction = "vssseg3e8.v,e64,m2";
	    34'b0100111???????101?01100110?????010  :  Instruction = "vssseg3e16.v,e64,m2";
	    34'b0100111???????110?01100110?????010  :  Instruction = "vssseg3e32.v,e64,m2";
	    34'b0100111???????111?01100110?????010  :  Instruction = "vssseg3e64.v,e64,m2";
	    34'b0100111???????000?01101010?????010  :  Instruction = "vssseg3e8.v,e64,m4";
	    34'b0100111???????101?01101010?????010  :  Instruction = "vssseg3e16.v,e64,m4";
	    34'b0100111???????110?01101010?????010  :  Instruction = "vssseg3e32.v,e64,m4";
	    34'b0100111???????000?01101110?????010  :  Instruction = "vssseg3e8.v,e64,m8";
	    34'b0100111???????101?01101110?????010  :  Instruction = "vssseg3e16.v,e64,m8";
	    34'b0100111???????111?011101?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e64,mf8";
	    34'b0100111???????110?011110?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e64,mf4";
	    34'b0100111???????111?011110?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e64,mf4";
	    34'b0100111???????101?011111?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e64,mf2";
	    34'b0100111???????110?011111?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e64,mf2";
	    34'b0100111???????111?011111?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e64,mf2";
	    34'b0100111???????000?011000?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e64,m1";
	    34'b0100111???????101?011000?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e64,m1";
	    34'b0100111???????110?011000?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e64,m1";
	    34'b0100111???????111?011000?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e64,m1";
	    34'b0100111???????000?011001?1?????010  :  Instruction = "vs[uo]xseg3ei8.v,e64,m2";
	    34'b0100111???????101?011001?1?????010  :  Instruction = "vs[uo]xseg3ei16.v,e64,m2";
	    34'b0100111???????110?011001?1?????010  :  Instruction = "vs[uo]xseg3ei32.v,e64,m2";
	    34'b0100111???????111?011001?1?????010  :  Instruction = "vs[uo]xseg3ei64.v,e64,m2";
	    34'b0100111???????111?01110100?0000011  :  Instruction = "vsseg4e64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000011  :  Instruction = "vsseg4e32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000011  :  Instruction = "vsseg4e64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000011  :  Instruction = "vsseg4e16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000011  :  Instruction = "vsseg4e32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000011  :  Instruction = "vsseg4e64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000011  :  Instruction = "vsseg4e8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000011  :  Instruction = "vsseg4e16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000011  :  Instruction = "vsseg4e32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000011  :  Instruction = "vsseg4e64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000011  :  Instruction = "vsseg4e8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000011  :  Instruction = "vsseg4e16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000011  :  Instruction = "vsseg4e32[ff].v,e64,m2";
	    34'b0100111???????111?01100100?0000011  :  Instruction = "vsseg4e64[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000011  :  Instruction = "vsseg4e8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000011  :  Instruction = "vsseg4e16[ff].v,e64,m4";
	    34'b0100111???????110?01101000?0000011  :  Instruction = "vsseg4e32[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000011  :  Instruction = "vsseg4e8[ff].v,e64,m8";
	    34'b0100111???????101?01101100?0000011  :  Instruction = "vsseg4e16[ff].v,e64,m8";
	    34'b0100111???????111?01110110?????011  :  Instruction = "vssseg4e64.v,e64,mf8";
	    34'b0100111???????110?01111010?????011  :  Instruction = "vssseg4e32.v,e64,mf4";
	    34'b0100111???????111?01111010?????011  :  Instruction = "vssseg4e64.v,e64,mf4";
	    34'b0100111???????101?01111110?????011  :  Instruction = "vssseg4e16.v,e64,mf2";
	    34'b0100111???????110?01111110?????011  :  Instruction = "vssseg4e32.v,e64,mf2";
	    34'b0100111???????111?01111110?????011  :  Instruction = "vssseg4e64.v,e64,mf2";
	    34'b0100111???????000?01100010?????011  :  Instruction = "vssseg4e8.v,e64,m1";
	    34'b0100111???????101?01100010?????011  :  Instruction = "vssseg4e16.v,e64,m1";
	    34'b0100111???????110?01100010?????011  :  Instruction = "vssseg4e32.v,e64,m1";
	    34'b0100111???????111?01100010?????011  :  Instruction = "vssseg4e64.v,e64,m1";
	    34'b0100111???????000?01100110?????011  :  Instruction = "vssseg4e8.v,e64,m2";
	    34'b0100111???????101?01100110?????011  :  Instruction = "vssseg4e16.v,e64,m2";
	    34'b0100111???????110?01100110?????011  :  Instruction = "vssseg4e32.v,e64,m2";
	    34'b0100111???????111?01100110?????011  :  Instruction = "vssseg4e64.v,e64,m2";
	    34'b0100111???????000?01101010?????011  :  Instruction = "vssseg4e8.v,e64,m4";
	    34'b0100111???????101?01101010?????011  :  Instruction = "vssseg4e16.v,e64,m4";
	    34'b0100111???????110?01101010?????011  :  Instruction = "vssseg4e32.v,e64,m4";
	    34'b0100111???????000?01101110?????011  :  Instruction = "vssseg4e8.v,e64,m8";
	    34'b0100111???????101?01101110?????011  :  Instruction = "vssseg4e16.v,e64,m8";
	    34'b0100111???????000?011???0001000011  :  Instruction = "vs4r.v,e64";
	    34'b0100111???????111?011101?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e64,mf8";
	    34'b0100111???????110?011110?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e64,mf4";
	    34'b0100111???????111?011110?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e64,mf4";
	    34'b0100111???????101?011111?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e64,mf2";
	    34'b0100111???????110?011111?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e64,mf2";
	    34'b0100111???????111?011111?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e64,mf2";
	    34'b0100111???????000?011000?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e64,m1";
	    34'b0100111???????101?011000?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e64,m1";
	    34'b0100111???????110?011000?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e64,m1";
	    34'b0100111???????111?011000?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e64,m1";
	    34'b0100111???????000?011001?1?????011  :  Instruction = "vs[uo]xseg4ei8.v,e64,m2";
	    34'b0100111???????101?011001?1?????011  :  Instruction = "vs[uo]xseg4ei16.v,e64,m2";
	    34'b0100111???????110?011001?1?????011  :  Instruction = "vs[uo]xseg4ei32.v,e64,m2";
	    34'b0100111???????111?011001?1?????011  :  Instruction = "vs[uo]xseg4ei64.v,e64,m2";
	    34'b0100111???????111?01110100?0000100  :  Instruction = "vsseg5e64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000100  :  Instruction = "vsseg5e32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000100  :  Instruction = "vsseg5e64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000100  :  Instruction = "vsseg5e16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000100  :  Instruction = "vsseg5e32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000100  :  Instruction = "vsseg5e64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000100  :  Instruction = "vsseg5e8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000100  :  Instruction = "vsseg5e16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000100  :  Instruction = "vsseg5e32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000100  :  Instruction = "vsseg5e64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000100  :  Instruction = "vsseg5e8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000100  :  Instruction = "vsseg5e16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000100  :  Instruction = "vsseg5e32[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000100  :  Instruction = "vsseg5e8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000100  :  Instruction = "vsseg5e16[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000100  :  Instruction = "vsseg5e8[ff].v,e64,m8";
	    34'b0100111???????111?01110110?????100  :  Instruction = "vssseg5e64.v,e64,mf8";
	    34'b0100111???????110?01111010?????100  :  Instruction = "vssseg5e32.v,e64,mf4";
	    34'b0100111???????111?01111010?????100  :  Instruction = "vssseg5e64.v,e64,mf4";
	    34'b0100111???????101?01111110?????100  :  Instruction = "vssseg5e16.v,e64,mf2";
	    34'b0100111???????110?01111110?????100  :  Instruction = "vssseg5e32.v,e64,mf2";
	    34'b0100111???????111?01111110?????100  :  Instruction = "vssseg5e64.v,e64,mf2";
	    34'b0100111???????000?01100010?????100  :  Instruction = "vssseg5e8.v,e64,m1";
	    34'b0100111???????101?01100010?????100  :  Instruction = "vssseg5e16.v,e64,m1";
	    34'b0100111???????110?01100010?????100  :  Instruction = "vssseg5e32.v,e64,m1";
	    34'b0100111???????111?01100010?????100  :  Instruction = "vssseg5e64.v,e64,m1";
	    34'b0100111???????000?01100110?????100  :  Instruction = "vssseg5e8.v,e64,m2";
	    34'b0100111???????101?01100110?????100  :  Instruction = "vssseg5e16.v,e64,m2";
	    34'b0100111???????110?01100110?????100  :  Instruction = "vssseg5e32.v,e64,m2";
	    34'b0100111???????000?01101010?????100  :  Instruction = "vssseg5e8.v,e64,m4";
	    34'b0100111???????101?01101010?????100  :  Instruction = "vssseg5e16.v,e64,m4";
	    34'b0100111???????000?01101110?????100  :  Instruction = "vssseg5e8.v,e64,m8";
	    34'b0100111???????111?011101?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e64,mf8";
	    34'b0100111???????110?011110?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e64,mf4";
	    34'b0100111???????111?011110?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e64,mf4";
	    34'b0100111???????101?011111?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e64,mf2";
	    34'b0100111???????110?011111?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e64,mf2";
	    34'b0100111???????111?011111?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e64,mf2";
	    34'b0100111???????000?011000?1?????100  :  Instruction = "vs[uo]xseg5ei8.v,e64,m1";
	    34'b0100111???????101?011000?1?????100  :  Instruction = "vs[uo]xseg5ei16.v,e64,m1";
	    34'b0100111???????110?011000?1?????100  :  Instruction = "vs[uo]xseg5ei32.v,e64,m1";
	    34'b0100111???????111?011000?1?????100  :  Instruction = "vs[uo]xseg5ei64.v,e64,m1";
	    34'b0100111???????111?01110100?0000101  :  Instruction = "vsseg6e64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000101  :  Instruction = "vsseg6e32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000101  :  Instruction = "vsseg6e64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000101  :  Instruction = "vsseg6e16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000101  :  Instruction = "vsseg6e32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000101  :  Instruction = "vsseg6e64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000101  :  Instruction = "vsseg6e8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000101  :  Instruction = "vsseg6e16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000101  :  Instruction = "vsseg6e32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000101  :  Instruction = "vsseg6e64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000101  :  Instruction = "vsseg6e8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000101  :  Instruction = "vsseg6e16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000101  :  Instruction = "vsseg6e32[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000101  :  Instruction = "vsseg6e8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000101  :  Instruction = "vsseg6e16[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000101  :  Instruction = "vsseg6e8[ff].v,e64,m8";
	    34'b0100111???????111?01110110?????101  :  Instruction = "vssseg6e64.v,e64,mf8";
	    34'b0100111???????110?01111010?????101  :  Instruction = "vssseg6e32.v,e64,mf4";
	    34'b0100111???????111?01111010?????101  :  Instruction = "vssseg6e64.v,e64,mf4";
	    34'b0100111???????101?01111110?????101  :  Instruction = "vssseg6e16.v,e64,mf2";
	    34'b0100111???????110?01111110?????101  :  Instruction = "vssseg6e32.v,e64,mf2";
	    34'b0100111???????111?01111110?????101  :  Instruction = "vssseg6e64.v,e64,mf2";
	    34'b0100111???????000?01100010?????101  :  Instruction = "vssseg6e8.v,e64,m1";
	    34'b0100111???????101?01100010?????101  :  Instruction = "vssseg6e16.v,e64,m1";
	    34'b0100111???????110?01100010?????101  :  Instruction = "vssseg6e32.v,e64,m1";
	    34'b0100111???????111?01100010?????101  :  Instruction = "vssseg6e64.v,e64,m1";
	    34'b0100111???????000?01100110?????101  :  Instruction = "vssseg6e8.v,e64,m2";
	    34'b0100111???????101?01100110?????101  :  Instruction = "vssseg6e16.v,e64,m2";
	    34'b0100111???????110?01100110?????101  :  Instruction = "vssseg6e32.v,e64,m2";
	    34'b0100111???????000?01101010?????101  :  Instruction = "vssseg6e8.v,e64,m4";
	    34'b0100111???????101?01101010?????101  :  Instruction = "vssseg6e16.v,e64,m4";
	    34'b0100111???????000?01101110?????101  :  Instruction = "vssseg6e8.v,e64,m8";
	    34'b0100111???????111?011101?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e64,mf8";
	    34'b0100111???????110?011110?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e64,mf4";
	    34'b0100111???????111?011110?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e64,mf4";
	    34'b0100111???????101?011111?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e64,mf2";
	    34'b0100111???????110?011111?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e64,mf2";
	    34'b0100111???????111?011111?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e64,mf2";
	    34'b0100111???????000?011000?1?????101  :  Instruction = "vs[uo]xseg6ei8.v,e64,m1";
	    34'b0100111???????101?011000?1?????101  :  Instruction = "vs[uo]xseg6ei16.v,e64,m1";
	    34'b0100111???????110?011000?1?????101  :  Instruction = "vs[uo]xseg6ei32.v,e64,m1";
	    34'b0100111???????111?011000?1?????101  :  Instruction = "vs[uo]xseg6ei64.v,e64,m1";
	    34'b0100111???????111?01110100?0000110  :  Instruction = "vsseg7e64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000110  :  Instruction = "vsseg7e32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000110  :  Instruction = "vsseg7e64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000110  :  Instruction = "vsseg7e16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000110  :  Instruction = "vsseg7e32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000110  :  Instruction = "vsseg7e64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000110  :  Instruction = "vsseg7e8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000110  :  Instruction = "vsseg7e16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000110  :  Instruction = "vsseg7e32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000110  :  Instruction = "vsseg7e64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000110  :  Instruction = "vsseg7e8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000110  :  Instruction = "vsseg7e16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000110  :  Instruction = "vsseg7e32[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000110  :  Instruction = "vsseg7e8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000110  :  Instruction = "vsseg7e16[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000110  :  Instruction = "vsseg7e8[ff].v,e64,m8";
	    34'b0100111???????111?01110110?????110  :  Instruction = "vssseg7e64.v,e64,mf8";
	    34'b0100111???????110?01111010?????110  :  Instruction = "vssseg7e32.v,e64,mf4";
	    34'b0100111???????111?01111010?????110  :  Instruction = "vssseg7e64.v,e64,mf4";
	    34'b0100111???????101?01111110?????110  :  Instruction = "vssseg7e16.v,e64,mf2";
	    34'b0100111???????110?01111110?????110  :  Instruction = "vssseg7e32.v,e64,mf2";
	    34'b0100111???????111?01111110?????110  :  Instruction = "vssseg7e64.v,e64,mf2";
	    34'b0100111???????000?01100010?????110  :  Instruction = "vssseg7e8.v,e64,m1";
	    34'b0100111???????101?01100010?????110  :  Instruction = "vssseg7e16.v,e64,m1";
	    34'b0100111???????110?01100010?????110  :  Instruction = "vssseg7e32.v,e64,m1";
	    34'b0100111???????111?01100010?????110  :  Instruction = "vssseg7e64.v,e64,m1";
	    34'b0100111???????000?01100110?????110  :  Instruction = "vssseg7e8.v,e64,m2";
	    34'b0100111???????101?01100110?????110  :  Instruction = "vssseg7e16.v,e64,m2";
	    34'b0100111???????110?01100110?????110  :  Instruction = "vssseg7e32.v,e64,m2";
	    34'b0100111???????000?01101010?????110  :  Instruction = "vssseg7e8.v,e64,m4";
	    34'b0100111???????101?01101010?????110  :  Instruction = "vssseg7e16.v,e64,m4";
	    34'b0100111???????000?01101110?????110  :  Instruction = "vssseg7e8.v,e64,m8";
	    34'b0100111???????111?011101?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e64,mf8";
	    34'b0100111???????110?011110?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e64,mf4";
	    34'b0100111???????111?011110?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e64,mf4";
	    34'b0100111???????101?011111?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e64,mf2";
	    34'b0100111???????110?011111?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e64,mf2";
	    34'b0100111???????111?011111?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e64,mf2";
	    34'b0100111???????000?011000?1?????110  :  Instruction = "vs[uo]xseg7ei8.v,e64,m1";
	    34'b0100111???????101?011000?1?????110  :  Instruction = "vs[uo]xseg7ei16.v,e64,m1";
	    34'b0100111???????110?011000?1?????110  :  Instruction = "vs[uo]xseg7ei32.v,e64,m1";
	    34'b0100111???????111?011000?1?????110  :  Instruction = "vs[uo]xseg7ei64.v,e64,m1";
	    34'b0100111???????111?01110100?0000111  :  Instruction = "vsseg8e64[ff].v,e64,mf8";
	    34'b0100111???????110?01111000?0000111  :  Instruction = "vsseg8e32[ff].v,e64,mf4";
	    34'b0100111???????111?01111000?0000111  :  Instruction = "vsseg8e64[ff].v,e64,mf4";
	    34'b0100111???????101?01111100?0000111  :  Instruction = "vsseg8e16[ff].v,e64,mf2";
	    34'b0100111???????110?01111100?0000111  :  Instruction = "vsseg8e32[ff].v,e64,mf2";
	    34'b0100111???????111?01111100?0000111  :  Instruction = "vsseg8e64[ff].v,e64,mf2";
	    34'b0100111???????000?01100000?0000111  :  Instruction = "vsseg8e8[ff].v,e64,m1";
	    34'b0100111???????101?01100000?0000111  :  Instruction = "vsseg8e16[ff].v,e64,m1";
	    34'b0100111???????110?01100000?0000111  :  Instruction = "vsseg8e32[ff].v,e64,m1";
	    34'b0100111???????111?01100000?0000111  :  Instruction = "vsseg8e64[ff].v,e64,m1";
	    34'b0100111???????000?01100100?0000111  :  Instruction = "vsseg8e8[ff].v,e64,m2";
	    34'b0100111???????101?01100100?0000111  :  Instruction = "vsseg8e16[ff].v,e64,m2";
	    34'b0100111???????110?01100100?0000111  :  Instruction = "vsseg8e32[ff].v,e64,m2";
	    34'b0100111???????000?01101000?0000111  :  Instruction = "vsseg8e8[ff].v,e64,m4";
	    34'b0100111???????101?01101000?0000111  :  Instruction = "vsseg8e16[ff].v,e64,m4";
	    34'b0100111???????000?01101100?0000111  :  Instruction = "vsseg8e8[ff].v,e64,m8";
	    34'b0100111???????000?011???0001000111  :  Instruction = "vs8r.v,e64";
	    34'b0100111???????111?01110110?????111  :  Instruction = "vssseg8e64.v,e64,mf8";
	    34'b0100111???????110?01111010?????111  :  Instruction = "vssseg8e32.v,e64,mf4";
	    34'b0100111???????111?01111010?????111  :  Instruction = "vssseg8e64.v,e64,mf4";
	    34'b0100111???????101?01111110?????111  :  Instruction = "vssseg8e16.v,e64,mf2";
	    34'b0100111???????110?01111110?????111  :  Instruction = "vssseg8e32.v,e64,mf2";
	    34'b0100111???????111?01111110?????111  :  Instruction = "vssseg8e64.v,e64,mf2";
	    34'b0100111???????000?01100010?????111  :  Instruction = "vssseg8e8.v,e64,m1";
	    34'b0100111???????101?01100010?????111  :  Instruction = "vssseg8e16.v,e64,m1";
	    34'b0100111???????110?01100010?????111  :  Instruction = "vssseg8e32.v,e64,m1";
	    34'b0100111???????111?01100010?????111  :  Instruction = "vssseg8e64.v,e64,m1";
	    34'b0100111???????000?01100110?????111  :  Instruction = "vssseg8e8.v,e64,m2";
	    34'b0100111???????101?01100110?????111  :  Instruction = "vssseg8e16.v,e64,m2";
	    34'b0100111???????110?01100110?????111  :  Instruction = "vssseg8e32.v,e64,m2";
	    34'b0100111???????000?01101010?????111  :  Instruction = "vssseg8e8.v,e64,m4";
	    34'b0100111???????101?01101010?????111  :  Instruction = "vssseg8e16.v,e64,m4";
	    34'b0100111???????000?01101110?????111  :  Instruction = "vssseg8e8.v,e64,m8";
	    34'b0100111???????111?011101?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e64,mf8";
	    34'b0100111???????110?011110?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e64,mf4";
	    34'b0100111???????111?011110?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e64,mf4";
	    34'b0100111???????101?011111?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e64,mf2";
	    34'b0100111???????110?011111?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e64,mf2";
	    34'b0100111???????111?011111?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e64,mf2";
	    34'b0100111???????000?011000?1?????111  :  Instruction = "vs[uo]xseg8ei8.v,e64,m1";
	    34'b0100111???????101?011000?1?????111  :  Instruction = "vs[uo]xseg8ei16.v,e64,m1";
	    34'b0100111???????110?011000?1?????111  :  Instruction = "vs[uo]xseg8ei32.v,e64,m1";
	    34'b0100111???????111?011000?1?????111  :  Instruction = "vs[uo]xseg8ei64.v,e64,m1";
	    default : Instruction = "ILLEG";
	endcase
end
//spyglass enable_block STARC05-2.10.3.2b_sa
//spyglass enable_block STARC05-2.10.3.2b_sb
//spyglass enable_block W164c
endmodule

module autogen_EncType (
input [6:0] Opcode,
input [2:0] funct3,
input [6:0] funct7,
input [1:0] mop,
output reg [4:0] EncType
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], mop[1], mop[0]})
	    18'b1010111010010000??  :  EncType[4] = 1'b1;
	    18'b1010111001010000??  :  EncType[4] = 1'b1;
	    18'b1010111?11100000??  :  EncType[4] = 1'b1;
	    18'b10101111?0010000??  :  EncType[4] = 1'b1;
	    18'b101011101101?111??  :  EncType[4] = 1'b1;
	    18'b101011110?10?111??  :  EncType[4] = 1'b1;
	    18'b10101110?00?0111??  :  EncType[4] = 1'b1;
	    18'b101011101100?011??  :  EncType[4] = 1'b1;
	    18'b101011110?01?111??  :  EncType[4] = 1'b1;
	    18'b0?00111000??????10  :  EncType[4] = 1'b1;
	    18'b1010111100?001?1??  :  EncType[4] = 1'b1;
	    18'b1010111010??1011??  :  EncType[4] = 1'b1;
	    18'b1010111011?00000??  :  EncType[4] = 1'b1;
	    18'b10101111011??100??  :  EncType[4] = 1'b1;
	    18'b10101110011??100??  :  EncType[4] = 1'b1;
	    18'b101011100111?1?0??  :  EncType[4] = 1'b1;
	    18'b1010111010??0100??  :  EncType[4] = 1'b1;
	    18'b1010111101110??0??  :  EncType[4] = 1'b1;
	    18'b10101110??001010??  :  EncType[4] = 1'b1;
	    18'b10101110011100????  :  EncType[4] = 1'b1;
	    18'b1010111010?11?00??  :  EncType[4] = 1'b1;
	    18'b1010111010?1?010??  :  EncType[4] = 1'b1;
	    18'b101011100?0110?1??  :  EncType[4] = 1'b1;
	    18'b101011100?01001???  :  EncType[4] = 1'b1;
	    18'b1010111101?11?00??  :  EncType[4] = 1'b1;
	    18'b1010111000?011?0??  :  EncType[4] = 1'b1;
	    18'b10101111000?11?0??  :  EncType[4] = 1'b1;
	    18'b1010111000?1000???  :  EncType[4] = 1'b1;
	    18'b1010111101?0100???  :  EncType[4] = 1'b1;
	    18'b1010111001??1000??  :  EncType[4] = 1'b1;
	    18'b101011110?01?000??  :  EncType[4] = 1'b1;
	    18'b101011101110?1?1??  :  EncType[4] = 1'b1;
	    18'b10101111100010????  :  EncType[4] = 1'b1;
	    18'b1010111000?000?0??  :  EncType[4] = 1'b1;
	    18'b0000111000??????00  :  EncType[4] = 1'b1;
	    18'b0?0011111???????10  :  EncType[4] = 1'b1;
	    18'b0100111000???????1  :  EncType[4] = 1'b1;
	    18'b10101111101??1?1??  :  EncType[4] = 1'b1;
	    18'b10101110101??1?1??  :  EncType[4] = 1'b1;
	    18'b0100111000???????0  :  EncType[4] = 1'b1;
	    18'b1010111011?011?0??  :  EncType[4] = 1'b1;
	    18'b101011101110?00???  :  EncType[4] = 1'b1;
	    18'b101011111011??1???  :  EncType[4] = 1'b1;
	    18'b101011110??0111???  :  EncType[4] = 1'b1;
	    18'b10101111101?01????  :  EncType[4] = 1'b1;
	    18'b10101110???01001??  :  EncType[4] = 1'b1;
	    18'b10101111011?11????  :  EncType[4] = 1'b1;
	    18'b101011100010???1??  :  EncType[4] = 1'b1;
	    18'b10101110011?11????  :  EncType[4] = 1'b1;
	    18'b1010111110110?????  :  EncType[4] = 1'b1;
	    18'b1010111010110?????  :  EncType[4] = 1'b1;
	    18'b1010111010?001????  :  EncType[4] = 1'b1;
	    18'b101011101101?00???  :  EncType[4] = 1'b1;
	    18'b10101111?0?010?1??  :  EncType[4] = 1'b1;
	    18'b101011110??01?10??  :  EncType[4] = 1'b1;
	    18'b101011110?011??1??  :  EncType[4] = 1'b1;
	    18'b101011101?0111????  :  EncType[4] = 1'b1;
	    18'b101011111111??????  :  EncType[4] = 1'b1;
	    18'b10101111?0001?1???  :  EncType[4] = 1'b1;
	    18'b101011111011???0??  :  EncType[4] = 1'b1;
	    18'b10101110?00001????  :  EncType[4] = 1'b1;
	    18'b10101110??011?00??  :  EncType[4] = 1'b1;
	    18'b10101110?0011?0???  :  EncType[4] = 1'b1;
	    18'b10101110?00?101???  :  EncType[4] = 1'b1;
	    18'b101011110010?0????  :  EncType[4] = 1'b1;
	    18'b101011110?000??0??  :  EncType[4] = 1'b1;
	    18'b10101111000??01???  :  EncType[4] = 1'b1;
	    18'b1010111001000?????  :  EncType[4] = 1'b1;
	    18'b0000111000???????1  :  EncType[4] = 1'b1;
	    18'b000011111???????00  :  EncType[4] = 1'b1;
	    18'b101011101000?0????  :  EncType[4] = 1'b1;
	    18'b010011111????????1  :  EncType[4] = 1'b1;
	    18'b101011110001?0????  :  EncType[4] = 1'b1;
	    18'b010011111????????0  :  EncType[4] = 1'b1;
	    18'b10101111110???????  :  EncType[4] = 1'b1;
	    18'b1010111011?01?1???  :  EncType[4] = 1'b1;
	    18'b101011110?101?????  :  EncType[4] = 1'b1;
	    18'b101011100?101?????  :  EncType[4] = 1'b1;
	    18'b000011111????????1  :  EncType[4] = 1'b1;
	    18'b0000000???????????  :  EncType[4] = 1'b1;
	    18'b0?001111?1????????  :  EncType[4] = 1'b1;
	    default : EncType[4] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], mop[0]})
	    18'b01100111?00100000?  :  EncType[3] = 1'b1;
	    18'b01100110??0000001?  :  EncType[3] = 1'b1;
	    18'b0110011?100010000?  :  EncType[3] = 1'b1;
	    18'b011001111?0100000?  :  EncType[3] = 1'b1;
	    18'b01100111??0000101?  :  EncType[3] = 1'b1;
	    18'b01100111?00010000?  :  EncType[3] = 1'b1;
	    18'b0110011100000010??  :  EncType[3] = 1'b1;
	    18'b0?10011?010110000?  :  EncType[3] = 1'b1;
	    18'b1010111010010000??  :  EncType[3] = 1'b1;
	    18'b1010111001010000??  :  EncType[3] = 1'b1;
	    18'b00100111010?101???  :  EncType[3] = 1'b1;
	    18'b00100111010110????  :  EncType[3] = 1'b1;
	    18'b10101111?0010000??  :  EncType[3] = 1'b1;
	    18'b101011101101?111??  :  EncType[3] = 1'b1;
	    18'b101011110?10?111??  :  EncType[3] = 1'b1;
	    18'b10101110?00?0111??  :  EncType[3] = 1'b1;
	    18'b101011101100?011??  :  EncType[3] = 1'b1;
	    18'b101011110?01?111??  :  EncType[3] = 1'b1;
	    18'b1010111100?001?1??  :  EncType[3] = 1'b1;
	    18'b1010111010??1011??  :  EncType[3] = 1'b1;
	    18'b1010111011?00000??  :  EncType[3] = 1'b1;
	    18'b10101111011??100??  :  EncType[3] = 1'b1;
	    18'b10101110011??100??  :  EncType[3] = 1'b1;
	    18'b101011100111?1?0??  :  EncType[3] = 1'b1;
	    18'b1010111010??0100??  :  EncType[3] = 1'b1;
	    18'b1010111101110??0??  :  EncType[3] = 1'b1;
	    18'b10101110??001010??  :  EncType[3] = 1'b1;
	    18'b10101110011100????  :  EncType[3] = 1'b1;
	    18'b1010111010?11?00??  :  EncType[3] = 1'b1;
	    18'b1010111010?1?010??  :  EncType[3] = 1'b1;
	    18'b101011100?0110?1??  :  EncType[3] = 1'b1;
	    18'b101011100?01001???  :  EncType[3] = 1'b1;
	    18'b1010111101?11?00??  :  EncType[3] = 1'b1;
	    18'b1010111000?011?0??  :  EncType[3] = 1'b1;
	    18'b10101111000?11?0??  :  EncType[3] = 1'b1;
	    18'b1010111000?1000???  :  EncType[3] = 1'b1;
	    18'b1010111101?0100???  :  EncType[3] = 1'b1;
	    18'b1010111001??1000??  :  EncType[3] = 1'b1;
	    18'b101011110?01?000??  :  EncType[3] = 1'b1;
	    18'b101011101110?1?1??  :  EncType[3] = 1'b1;
	    18'b10101111100010????  :  EncType[3] = 1'b1;
	    18'b1010111000?000?0??  :  EncType[3] = 1'b1;
	    18'b0100111000???????1  :  EncType[3] = 1'b1;
	    18'b010?1111?1???????1  :  EncType[3] = 1'b1;
	    18'b10101111101??1?1??  :  EncType[3] = 1'b1;
	    18'b10101110101??1?1??  :  EncType[3] = 1'b1;
	    18'b1010111011?011?0??  :  EncType[3] = 1'b1;
	    18'b101011101110?00???  :  EncType[3] = 1'b1;
	    18'b101011111011??1???  :  EncType[3] = 1'b1;
	    18'b101011110??0111???  :  EncType[3] = 1'b1;
	    18'b10101111101?01????  :  EncType[3] = 1'b1;
	    18'b10101110???01001??  :  EncType[3] = 1'b1;
	    18'b10101111011?11????  :  EncType[3] = 1'b1;
	    18'b101011100010???1??  :  EncType[3] = 1'b1;
	    18'b10101110011?11????  :  EncType[3] = 1'b1;
	    18'b1010111110110?????  :  EncType[3] = 1'b1;
	    18'b1010111010110?????  :  EncType[3] = 1'b1;
	    18'b1010111010?001????  :  EncType[3] = 1'b1;
	    18'b101011101101?00???  :  EncType[3] = 1'b1;
	    18'b10101111?0?010?1??  :  EncType[3] = 1'b1;
	    18'b101011110??01?10??  :  EncType[3] = 1'b1;
	    18'b101011110?011??1??  :  EncType[3] = 1'b1;
	    18'b101011101?0111????  :  EncType[3] = 1'b1;
	    18'b10101111?0001?1???  :  EncType[3] = 1'b1;
	    18'b101011111011???0??  :  EncType[3] = 1'b1;
	    18'b10101110?00001????  :  EncType[3] = 1'b1;
	    18'b10101110??011?00??  :  EncType[3] = 1'b1;
	    18'b10101110?0011?0???  :  EncType[3] = 1'b1;
	    18'b10101110?00?101???  :  EncType[3] = 1'b1;
	    18'b101011110010?0????  :  EncType[3] = 1'b1;
	    18'b101011110?000??0??  :  EncType[3] = 1'b1;
	    18'b10101111000??01???  :  EncType[3] = 1'b1;
	    18'b1010111001000?????  :  EncType[3] = 1'b1;
	    18'b101011101000?0????  :  EncType[3] = 1'b1;
	    18'b010011111????????1  :  EncType[3] = 1'b1;
	    18'b101011110001?0????  :  EncType[3] = 1'b1;
	    18'b1010111011?01?1???  :  EncType[3] = 1'b1;
	    18'b101011110?101?????  :  EncType[3] = 1'b1;
	    18'b101011100?101?????  :  EncType[3] = 1'b1;
	    18'b0000000???????????  :  EncType[3] = 1'b1;
	    18'b0?00111010????????  :  EncType[3] = 1'b1;
	    18'b0?00111001????????  :  EncType[3] = 1'b1;
	    18'b0101111???????????  :  EncType[3] = 1'b1;
	    18'b10?0011???????????  :  EncType[3] = 1'b1;
	    18'b100??11???????????  :  EncType[3] = 1'b1;
	    default : EncType[3] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], mop[1], mop[0]})
	    18'b1010111010010000??  :  EncType[2] = 1'b1;
	    18'b1010111001010000??  :  EncType[2] = 1'b1;
	    18'b0?00111000??????10  :  EncType[2] = 1'b1;
	    18'b0?0011111???????10  :  EncType[2] = 1'b1;
	    18'b01001111?1???????0  :  EncType[2] = 1'b1;
	    18'b0100111000???????0  :  EncType[2] = 1'b1;
	    18'b0000111000???????1  :  EncType[2] = 1'b1;
	    18'b?0001111?1??????1?  :  EncType[2] = 1'b1;
	    18'b010011111????????0  :  EncType[2] = 1'b1;
	    18'b?0001111?1???????1  :  EncType[2] = 1'b1;
	    18'b000011111????????1  :  EncType[2] = 1'b1;
	    18'b0000000???????????  :  EncType[2] = 1'b1;
	    18'b0?00111010????????  :  EncType[2] = 1'b1;
	    18'b0?00111001????????  :  EncType[2] = 1'b1;
	    18'b1?01111???????????  :  EncType[2] = 1'b1;
	    18'b1?00011???????????  :  EncType[2] = 1'b1;
	    18'b0001111???????????  :  EncType[2] = 1'b1;
	    18'b10?0011???????????  :  EncType[2] = 1'b1;
	    18'b0?10111???????????  :  EncType[2] = 1'b1;
	    18'b100??11???????????  :  EncType[2] = 1'b1;
	    default : EncType[2] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], mop[1], mop[0]})
	    19'b01100111?00100000??  :  EncType[1] = 1'b1;
	    19'b0110011?100010000??  :  EncType[1] = 1'b1;
	    19'b011001111?0100000??  :  EncType[1] = 1'b1;
	    19'b01100111??0000101??  :  EncType[1] = 1'b1;
	    19'b01100111?00010000??  :  EncType[1] = 1'b1;
	    19'b0110011100000010???  :  EncType[1] = 1'b1;
	    19'b0?10011?010110000??  :  EncType[1] = 1'b1;
	    19'b10101??0010100?0???  :  EncType[1] = 1'b1;
	    19'b00?00?????0000000??  :  EncType[1] = 1'b1;
	    19'b00?00??1??0?00000??  :  EncType[1] = 1'b1;
	    19'b1010111?11100000???  :  EncType[1] = 1'b1;
	    19'b00100111010?101????  :  EncType[1] = 1'b1;
	    19'b10101??011?010?1???  :  EncType[1] = 1'b1;
	    19'b10101??0110111?????  :  EncType[1] = 1'b1;
	    19'b00100111010110?????  :  EncType[1] = 1'b1;
	    19'b10101111?0010000???  :  EncType[1] = 1'b1;
	    19'b101011101101?111???  :  EncType[1] = 1'b1;
	    19'b101011110?10?111???  :  EncType[1] = 1'b1;
	    19'b101011101100?011???  :  EncType[1] = 1'b1;
	    19'b101011110?01?111???  :  EncType[1] = 1'b1;
	    19'b1010111100?001?1???  :  EncType[1] = 1'b1;
	    19'b1010111011?00000???  :  EncType[1] = 1'b1;
	    19'b10101111011??100???  :  EncType[1] = 1'b1;
	    19'b1010111101110??0???  :  EncType[1] = 1'b1;
	    19'b1010111101?11?00???  :  EncType[1] = 1'b1;
	    19'b10101111000?11?0???  :  EncType[1] = 1'b1;
	    19'b1010111101?0100????  :  EncType[1] = 1'b1;
	    19'b101011110?01?000???  :  EncType[1] = 1'b1;
	    19'b101011101110?1?1???  :  EncType[1] = 1'b1;
	    19'b10101111100010?????  :  EncType[1] = 1'b1;
	    19'b0000111000???????00  :  EncType[1] = 1'b1;
	    19'b01001111?1????????0  :  EncType[1] = 1'b1;
	    19'b10101111101??1?1???  :  EncType[1] = 1'b1;
	    19'b0100111000????????0  :  EncType[1] = 1'b1;
	    19'b1010111011?011?0???  :  EncType[1] = 1'b1;
	    19'b101011101110?00????  :  EncType[1] = 1'b1;
	    19'b101011111011??1????  :  EncType[1] = 1'b1;
	    19'b101011110??0111????  :  EncType[1] = 1'b1;
	    19'b10101111101?01?????  :  EncType[1] = 1'b1;
	    19'b10101111011?11?????  :  EncType[1] = 1'b1;
	    19'b000?1??1?1???????00  :  EncType[1] = 1'b1;
	    19'b1010111110110??????  :  EncType[1] = 1'b1;
	    19'b101011101101?00????  :  EncType[1] = 1'b1;
	    19'b10101111?0?010?1???  :  EncType[1] = 1'b1;
	    19'b101011110??01?10???  :  EncType[1] = 1'b1;
	    19'b101011110?011??1???  :  EncType[1] = 1'b1;
	    19'b10101111?0001?1????  :  EncType[1] = 1'b1;
	    19'b101011111011???0???  :  EncType[1] = 1'b1;
	    19'b101011110010?0?????  :  EncType[1] = 1'b1;
	    19'b101011110?000??0???  :  EncType[1] = 1'b1;
	    19'b10101111000??01????  :  EncType[1] = 1'b1;
	    19'b000011111????????00  :  EncType[1] = 1'b1;
	    19'b101011110001?0?????  :  EncType[1] = 1'b1;
	    19'b010011111?????????0  :  EncType[1] = 1'b1;
	    19'b1010111011?01?1????  :  EncType[1] = 1'b1;
	    19'b101011110?101??????  :  EncType[1] = 1'b1;
	    19'b0?00111010?????????  :  EncType[1] = 1'b1;
	    19'b0?00111001?????????  :  EncType[1] = 1'b1;
	    19'b00?00???1??????????  :  EncType[1] = 1'b1;
	    19'b0001111????????????  :  EncType[1] = 1'b1;
	    19'b00?00????0?????????  :  EncType[1] = 1'b1;
	    19'b0?000??????????????  :  EncType[1] = 1'b1;
	    19'b110?1??????????????  :  EncType[1] = 1'b1;
	    19'b??????0????????????  :  EncType[1] = 1'b1;
	    19'b?????0?????????????  :  EncType[1] = 1'b1;
	    default : EncType[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], mop[1], mop[0]})
	    19'b01?00???010110000??  :  EncType[0] = 1'b1;
	    19'b01?00??10101?0000??  :  EncType[0] = 1'b1;
	    19'b0110011?100010000??  :  EncType[0] = 1'b1;
	    19'b011001111?0100000??  :  EncType[0] = 1'b1;
	    19'b01100111?00010000??  :  EncType[0] = 1'b1;
	    19'b01?00???000?00000??  :  EncType[0] = 1'b1;
	    19'b0110011100000010???  :  EncType[0] = 1'b1;
	    19'b01?00?????0000000??  :  EncType[0] = 1'b1;
	    19'b01?00??1??0000?01??  :  EncType[0] = 1'b1;
	    19'b010?1??1?1???????10  :  EncType[0] = 1'b1;
	    19'b010?1??11????????10  :  EncType[0] = 1'b1;
	    19'b101011101101?111???  :  EncType[0] = 1'b1;
	    19'b10101110?00?0111???  :  EncType[0] = 1'b1;
	    19'b101011101100?011???  :  EncType[0] = 1'b1;
	    19'b0100???00????????10  :  EncType[0] = 1'b1;
	    19'b1010111010??1011???  :  EncType[0] = 1'b1;
	    19'b1010111011?00000???  :  EncType[0] = 1'b1;
	    19'b10101110011??100???  :  EncType[0] = 1'b1;
	    19'b101011100111?1?0???  :  EncType[0] = 1'b1;
	    19'b1010111010??0100???  :  EncType[0] = 1'b1;
	    19'b10101110??001010???  :  EncType[0] = 1'b1;
	    19'b10101110011100?????  :  EncType[0] = 1'b1;
	    19'b1010111010?11?00???  :  EncType[0] = 1'b1;
	    19'b1010111010?1?010???  :  EncType[0] = 1'b1;
	    19'b101011100?0110?1???  :  EncType[0] = 1'b1;
	    19'b101011100?01001????  :  EncType[0] = 1'b1;
	    19'b1010111000?011?0???  :  EncType[0] = 1'b1;
	    19'b1010111000?1000????  :  EncType[0] = 1'b1;
	    19'b1010111001??1000???  :  EncType[0] = 1'b1;
	    19'b101011101110?1?1???  :  EncType[0] = 1'b1;
	    19'b1010111000?000?0???  :  EncType[0] = 1'b1;
	    19'b0000111000???????00  :  EncType[0] = 1'b1;
	    19'b10101110101??1?1???  :  EncType[0] = 1'b1;
	    19'b1010111011?011?0???  :  EncType[0] = 1'b1;
	    19'b010?1??010?????????  :  EncType[0] = 1'b1;
	    19'b101011101110?00????  :  EncType[0] = 1'b1;
	    19'b010?1??001?????????  :  EncType[0] = 1'b1;
	    19'b10101110???01001???  :  EncType[0] = 1'b1;
	    19'b000?1??1?1???????00  :  EncType[0] = 1'b1;
	    19'b101011100010???1???  :  EncType[0] = 1'b1;
	    19'b10101110011?11?????  :  EncType[0] = 1'b1;
	    19'b1010111010110??????  :  EncType[0] = 1'b1;
	    19'b1010111010?001?????  :  EncType[0] = 1'b1;
	    19'b101011101101?00????  :  EncType[0] = 1'b1;
	    19'b101011101?0111?????  :  EncType[0] = 1'b1;
	    19'b101011111111???????  :  EncType[0] = 1'b1;
	    19'b10101110?00001?????  :  EncType[0] = 1'b1;
	    19'b10101110??011?00???  :  EncType[0] = 1'b1;
	    19'b10101110?0011?0????  :  EncType[0] = 1'b1;
	    19'b10101110?00?101????  :  EncType[0] = 1'b1;
	    19'b1010111001000??????  :  EncType[0] = 1'b1;
	    19'b0000111000????????1  :  EncType[0] = 1'b1;
	    19'b000011111????????00  :  EncType[0] = 1'b1;
	    19'b101011101000?0?????  :  EncType[0] = 1'b1;
	    19'b1010111011?01?1????  :  EncType[0] = 1'b1;
	    19'b101011100?101??????  :  EncType[0] = 1'b1;
	    19'b?0001111?1????????1  :  EncType[0] = 1'b1;
	    19'b000011111?????????1  :  EncType[0] = 1'b1;
	    19'b01000??????????????  :  EncType[0] = 1'b1;
	    19'b0101111????????????  :  EncType[0] = 1'b1;
	    19'b0001111????????????  :  EncType[0] = 1'b1;
	    19'b0?10111????????????  :  EncType[0] = 1'b1;
	    19'b100??11????????????  :  EncType[0] = 1'b1;
	    19'b??????0????????????  :  EncType[0] = 1'b1;
	    19'b?????0?????????????  :  EncType[0] = 1'b1;
	    default : EncType[0] = 1'b0;
	endcase
end
endmodule

module autogen_SrcA (
input [6:0] Opcode,
input [2:0] funct3,
input [6:0] funct7,
output reg [1:0] SrcA
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0]})
	    17'b10?011110110?111?  :  SrcA[1] = 1'b1;
	    17'b10?01110?00?101??  :  SrcA[1] = 1'b1;
	    17'b10?011110101?111?  :  SrcA[1] = 1'b1;
	    17'b10?0111010?11?11?  :  SrcA[1] = 1'b1;
	    17'b10?0111101?0111??  :  SrcA[1] = 1'b1;
	    17'b10?01110?00?0111?  :  SrcA[1] = 1'b1;
	    17'b10?0111101?1110??  :  SrcA[1] = 1'b1;
	    17'b10?0111010?1110??  :  SrcA[1] = 1'b1;
	    17'b10?0111010?110?0?  :  SrcA[1] = 1'b1;
	    17'b10?0111?01101????  :  SrcA[1] = 1'b1;
	    17'b10?0111001000????  :  SrcA[1] = 1'b1;
	    17'b10?0111000?1000??  :  SrcA[1] = 1'b1;
	    17'b10?01110?0011?0??  :  SrcA[1] = 1'b1;
	    17'b10?0111101?1?000?  :  SrcA[1] = 1'b1;
	    17'b10?0111?011??100?  :  SrcA[1] = 1'b1;
	    17'b10?0011????1000?0  :  SrcA[1] = 1'b1;
	    17'b10?0111?01110??0?  :  SrcA[1] = 1'b1;
	    17'b10?0011???1?100?0  :  SrcA[1] = 1'b1;
	    17'b10?0111?01?0100??  :  SrcA[1] = 1'b1;
	    17'b10?011100?0001???  :  SrcA[1] = 1'b1;
	    17'b10?01110?0000??0?  :  SrcA[1] = 1'b1;
	    17'b10?0111?010110?1?  :  SrcA[1] = 1'b1;
	    17'b10?0111?01?11?00?  :  SrcA[1] = 1'b1;
	    17'b10?0111000?011?0?  :  SrcA[1] = 1'b1;
	    17'b10?01110011100???  :  SrcA[1] = 1'b1;
	    17'b10?0111010?001???  :  SrcA[1] = 1'b1;
	    17'b10?011101000?0???  :  SrcA[1] = 1'b1;
	    17'b10?0111010110????  :  SrcA[1] = 1'b1;
	    17'b10?0111?01000??0?  :  SrcA[1] = 1'b1;
	    17'b10?01110?010?1?1?  :  SrcA[1] = 1'b1;
	    17'b10?0111010011????  :  SrcA[1] = 1'b1;
	    17'b10?01110?0?010?1?  :  SrcA[1] = 1'b1;
	    17'b10?0111?01?010?0?  :  SrcA[1] = 1'b1;
	    17'b10?011100010?0???  :  SrcA[1] = 1'b1;
	    17'b10?011100001?0???  :  SrcA[1] = 1'b1;
	    17'b10?0111?011?11???  :  SrcA[1] = 1'b1;
	    17'b10?0011???00?0??0  :  SrcA[1] = 1'b1;
	    17'b10?0011???000?0?0  :  SrcA[1] = 1'b1;
	    17'b100??11??????????  :  SrcA[1] = 1'b1;
	    default : SrcA[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[3], funct7[2], funct7[0]})
	    15'b?0100?????11100  :  SrcA[0] = 1'b1;
	    15'b0?0?1??????????  :  SrcA[0] = 1'b1;
	    15'b?1?00??01??????  :  SrcA[0] = 1'b1;
	    15'b0??00??????????  :  SrcA[0] = 1'b1;
	    15'b?1?00??0?1?????  :  SrcA[0] = 1'b1;
	    15'b?100???????????  :  SrcA[0] = 1'b1;
	    15'b??????0????????  :  SrcA[0] = 1'b1;
	    15'b?????0?????????  :  SrcA[0] = 1'b1;
	    15'b10101??????????  :  SrcA[0] = 1'b1;
	    default : SrcA[0] = 1'b0;
	endcase
end
endmodule

module autogen_SrcB (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [1:0] mop,
input [0:0] vm,
output reg [1:0] SrcB
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0], mop[0], vm[0]})
	    19'b1010111??0111?010??  :  SrcB[1] = 1'b1;
	    19'b101011101?111?01??0  :  SrcB[1] = 1'b1;
	    19'b101011110?111?10???  :  SrcB[1] = 1'b1;
	    19'b10101110?0111??00?0  :  SrcB[1] = 1'b1;
	    19'b101011111??11??10??  :  SrcB[1] = 1'b1;
	    19'b10101110010????10??  :  SrcB[1] = 1'b1;
	    19'b10101110??01??100??  :  SrcB[1] = 1'b1;
	    19'b101011100?011?01???  :  SrcB[1] = 1'b1;
	    19'b10101111??100??01??  :  SrcB[1] = 1'b1;
	    19'b1010111?011?0?011??  :  SrcB[1] = 1'b1;
	    19'b101011101?111?101??  :  SrcB[1] = 1'b1;
	    19'b10101110?1?1??100??  :  SrcB[1] = 1'b1;
	    19'b10101110110?1??0???  :  SrcB[1] = 1'b1;
	    19'b1010111011?0???00??  :  SrcB[1] = 1'b1;
	    19'b101011111???0?110??  :  SrcB[1] = 1'b1;
	    19'b10101110?0000?0????  :  SrcB[1] = 1'b1;
	    19'b101011110?00??011??  :  SrcB[1] = 1'b1;
	    19'b101011110?1?1?01???  :  SrcB[1] = 1'b1;
	    19'b101011111000??00???  :  SrcB[1] = 1'b1;
	    19'b1010111001?1??1?0??  :  SrcB[1] = 1'b1;
	    19'b101011101?00??011??  :  SrcB[1] = 1'b1;
	    19'b1010111?0111??10???  :  SrcB[1] = 1'b1;
	    19'b1010111?1001??001??  :  SrcB[1] = 1'b1;
	    19'b1010111?1101??010??  :  SrcB[1] = 1'b1;
	    19'b1010111000????001??  :  SrcB[1] = 1'b1;
	    19'b1010111?1??00?010??  :  SrcB[1] = 1'b1;
	    19'b1010111110??0??01??  :  SrcB[1] = 1'b1;
	    19'b10101111??1?1??10??  :  SrcB[1] = 1'b1;
	    19'b1010111?11?00??01??  :  SrcB[1] = 1'b1;
	    19'b1010111110?????10??  :  SrcB[1] = 1'b1;
	    19'b1010111011?0??10???  :  SrcB[1] = 1'b1;
	    19'b10101110?1001?0????  :  SrcB[1] = 1'b1;
	    19'b10101110??0?0?010??  :  SrcB[1] = 1'b1;
	    19'b1010111?01010??0???  :  SrcB[1] = 1'b1;
	    19'b1010111?001?1??00??  :  SrcB[1] = 1'b1;
	    19'b1010111?01?1??011??  :  SrcB[1] = 1'b1;
	    19'b1010111?011?0??00??  :  SrcB[1] = 1'b1;
	    19'b1010111?0100???01??  :  SrcB[1] = 1'b1;
	    19'b1010111000????010??  :  SrcB[1] = 1'b1;
	    19'b10101110111???01???  :  SrcB[1] = 1'b1;
	    19'b10101111?01????10??  :  SrcB[1] = 1'b1;
	    19'b10101111?11????01??  :  SrcB[1] = 1'b1;
	    19'b1010111000??0??0???  :  SrcB[1] = 1'b1;
	    19'b1010111101?????0???  :  SrcB[1] = 1'b1;
	    19'b1010111?010?1???0??  :  SrcB[1] = 1'b1;
	    19'b101011110?0????00??  :  SrcB[1] = 1'b1;
	    19'b101011101?0????00??  :  SrcB[1] = 1'b1;
	    19'b10?0011000?0?0?????  :  SrcB[1] = 1'b1;
	    19'b10?001100?0??0?????  :  SrcB[1] = 1'b1;
	    19'b10?0011?0100?0?????  :  SrcB[1] = 1'b1;
	    19'b0100111???????010??  :  SrcB[1] = 1'b1;
	    19'b0?00111??????????1?  :  SrcB[1] = 1'b1;
	    19'b100??11????????????  :  SrcB[1] = 1'b1;
	    default : SrcB[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], mop[1], mop[0], vm[0]})
	    19'b010?1????????001???  :  SrcB[0] = 1'b1;
	    19'b1010111??0111010???  :  SrcB[0] = 1'b1;
	    19'b101011101?11101???0  :  SrcB[0] = 1'b1;
	    19'b101011110?11110????  :  SrcB[0] = 1'b1;
	    19'b10101110?0111?00??0  :  SrcB[0] = 1'b1;
	    19'b101011111??11?10???  :  SrcB[0] = 1'b1;
	    19'b10101110010???10???  :  SrcB[0] = 1'b1;
	    19'b10101110??01?100???  :  SrcB[0] = 1'b1;
	    19'b101011100?01101????  :  SrcB[0] = 1'b1;
	    19'b10101111??100?01???  :  SrcB[0] = 1'b1;
	    19'b1010111?011?0011???  :  SrcB[0] = 1'b1;
	    19'b101011101?111101???  :  SrcB[0] = 1'b1;
	    19'b10101110?1?1?100???  :  SrcB[0] = 1'b1;
	    19'b10101110110?1?0????  :  SrcB[0] = 1'b1;
	    19'b1010111011?0??00???  :  SrcB[0] = 1'b1;
	    19'b101011111???0110???  :  SrcB[0] = 1'b1;
	    19'b10101110?00000?????  :  SrcB[0] = 1'b1;
	    19'b101011110?00?011???  :  SrcB[0] = 1'b1;
	    19'b101011110?1?101????  :  SrcB[0] = 1'b1;
	    19'b101011111000?00????  :  SrcB[0] = 1'b1;
	    19'b1010111001?1?1?0???  :  SrcB[0] = 1'b1;
	    19'b101011101?00?011???  :  SrcB[0] = 1'b1;
	    19'b1010111?0111?10????  :  SrcB[0] = 1'b1;
	    19'b1010111?1001?001???  :  SrcB[0] = 1'b1;
	    19'b1010111?1101?010???  :  SrcB[0] = 1'b1;
	    19'b1010111000???001???  :  SrcB[0] = 1'b1;
	    19'b1010111?1??00010???  :  SrcB[0] = 1'b1;
	    19'b1010111110??0?01???  :  SrcB[0] = 1'b1;
	    19'b10101111??1?1?10???  :  SrcB[0] = 1'b1;
	    19'b1010111?11?00?01???  :  SrcB[0] = 1'b1;
	    19'b1010111110????10???  :  SrcB[0] = 1'b1;
	    19'b1010111011?0?10????  :  SrcB[0] = 1'b1;
	    19'b10101110?10010?????  :  SrcB[0] = 1'b1;
	    19'b10101110??0?0010???  :  SrcB[0] = 1'b1;
	    19'b1010111?01010?0????  :  SrcB[0] = 1'b1;
	    19'b1010111?001?1?00???  :  SrcB[0] = 1'b1;
	    19'b1010111?01?1?011???  :  SrcB[0] = 1'b1;
	    19'b1010111?011?0?00???  :  SrcB[0] = 1'b1;
	    19'b1010111?0100??01???  :  SrcB[0] = 1'b1;
	    19'b1010111000???010???  :  SrcB[0] = 1'b1;
	    19'b10101110111??01????  :  SrcB[0] = 1'b1;
	    19'b10101111?01???10???  :  SrcB[0] = 1'b1;
	    19'b10101111?11???01???  :  SrcB[0] = 1'b1;
	    19'b1010111000??0?0????  :  SrcB[0] = 1'b1;
	    19'b1010111101????0????  :  SrcB[0] = 1'b1;
	    19'b1010111?010?1??0???  :  SrcB[0] = 1'b1;
	    19'b101011110?0???00???  :  SrcB[0] = 1'b1;
	    19'b101011101?0???00???  :  SrcB[0] = 1'b1;
	    19'b10101??100000?11???  :  SrcB[0] = 1'b1;
	    19'b0?001???????????1??  :  SrcB[0] = 1'b1;
	    19'b0?00111??????????1?  :  SrcB[0] = 1'b1;
	    19'b01011??????????????  :  SrcB[0] = 1'b1;
	    19'b01?00??????????????  :  SrcB[0] = 1'b1;
	    19'b?1000??????????????  :  SrcB[0] = 1'b1;
	    19'b??????0????????????  :  SrcB[0] = 1'b1;
	    19'b?????0?????????????  :  SrcB[0] = 1'b1;
	    default : SrcB[0] = 1'b0;
	endcase
end
endmodule

module autogen_SrcC (
input [6:0] Opcode,
input [2:0] funct3,
output reg [1:0] SrcC
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0]})
	    10'b0100111000  :  SrcC[1] = 1'b1;
	    10'b010011111?  :  SrcC[1] = 1'b1;
	    10'b01001111?1  :  SrcC[1] = 1'b1;
	    10'b100??11???  :  SrcC[1] = 1'b1;
	    default : SrcC[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0]})
	    10'b0100111000  :  SrcC[0] = 1'b1;
	    10'b010011111?  :  SrcC[0] = 1'b1;
	    10'b01001111?1  :  SrcC[0] = 1'b1;
	    default : SrcC[0] = 1'b0;
	endcase
end
endmodule

module autogen_Dest (
input [6:0] Opcode,
input [2:0] funct3,
input [6:0] funct7,
output reg [1:0] Dest
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0]})
	    17'b10?0111010??0100?  :  Dest[1] = 1'b1;
	    17'b101011110?10?111?  :  Dest[1] = 1'b1;
	    17'b1010111?1011??11?  :  Dest[1] = 1'b1;
	    17'b101011110?01?000?  :  Dest[1] = 1'b1;
	    17'b101011101?00?011?  :  Dest[1] = 1'b1;
	    17'b10101111?0010000?  :  Dest[1] = 1'b1;
	    17'b1010111?000?0111?  :  Dest[1] = 1'b1;
	    17'b10?01110?10?0000?  :  Dest[1] = 1'b1;
	    17'b1010111?011??100?  :  Dest[1] = 1'b1;
	    17'b10?0111010?11?00?  :  Dest[1] = 1'b1;
	    17'b101011101?01?111?  :  Dest[1] = 1'b1;
	    17'b101011110??0111??  :  Dest[1] = 1'b1;
	    17'b1010111011?011?0?  :  Dest[1] = 1'b1;
	    17'b10101111000?1?1??  :  Dest[1] = 1'b1;
	    17'b1010111?0?0110?1?  :  Dest[1] = 1'b1;
	    17'b1010111?100010???  :  Dest[1] = 1'b1;
	    17'b101011110?01?111?  :  Dest[1] = 1'b1;
	    17'b101011101?10?1?1?  :  Dest[1] = 1'b1;
	    17'b101011111011???0?  :  Dest[1] = 1'b1;
	    17'b10101111000???11?  :  Dest[1] = 1'b1;
	    17'b101011101110?00??  :  Dest[1] = 1'b1;
	    17'b101011110?011??1?  :  Dest[1] = 1'b1;
	    17'b101011100?11000??  :  Dest[1] = 1'b1;
	    17'b1010111?0??01010?  :  Dest[1] = 1'b1;
	    17'b1010111001000????  :  Dest[1] = 1'b1;
	    17'b1010111001?1001??  :  Dest[1] = 1'b1;
	    17'b101011101101?00??  :  Dest[1] = 1'b1;
	    17'b1010111010?1101??  :  Dest[1] = 1'b1;
	    17'b1010111?101?01???  :  Dest[1] = 1'b1;
	    17'b10101111?0001?1??  :  Dest[1] = 1'b1;
	    17'b1010111?01110??0?  :  Dest[1] = 1'b1;
	    17'b1010111?00?001?1?  :  Dest[1] = 1'b1;
	    17'b10101110??0?1001?  :  Dest[1] = 1'b1;
	    17'b1010111011?01?1??  :  Dest[1] = 1'b1;
	    17'b1010111?10110????  :  Dest[1] = 1'b1;
	    17'b?000111?10???????  :  Dest[1] = 1'b1;
	    17'b1010111?01?11?00?  :  Dest[1] = 1'b1;
	    17'b10101110?00??010?  :  Dest[1] = 1'b1;
	    17'b101011101?0111???  :  Dest[1] = 1'b1;
	    17'b?00011100????????  :  Dest[1] = 1'b1;
	    17'b1010111?00?011?0?  :  Dest[1] = 1'b1;
	    17'b1010111?01?0100??  :  Dest[1] = 1'b1;
	    17'b1010111010000????  :  Dest[1] = 1'b1;
	    17'b1010111?00011?0??  :  Dest[1] = 1'b1;
	    17'b1010111?0001?0???  :  Dest[1] = 1'b1;
	    17'b1010111?101??1?1?  :  Dest[1] = 1'b1;
	    17'b1010111?011?11???  :  Dest[1] = 1'b1;
	    17'b1010111?0?101????  :  Dest[1] = 1'b1;
	    17'b1010111??0?010?1?  :  Dest[1] = 1'b1;
	    17'b00001111?1???????  :  Dest[1] = 1'b1;
	    17'b1010111?0?000??0?  :  Dest[1] = 1'b1;
	    17'b1010111?0010?0???  :  Dest[1] = 1'b1;
	    17'b10?0011???11?10?0  :  Dest[1] = 1'b1;
	    17'b10?0011???0?000?0  :  Dest[1] = 1'b1;
	    17'b10?0011???000?0?0  :  Dest[1] = 1'b1;
	    17'b10?0011???00?0??0  :  Dest[1] = 1'b1;
	    17'b100??11??????????  :  Dest[1] = 1'b1;
	    default : Dest[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0]})
	    17'b101011110?10?111?  :  Dest[0] = 1'b1;
	    17'b?010011???1?100?0  :  Dest[0] = 1'b1;
	    17'b1010111?1011??11?  :  Dest[0] = 1'b1;
	    17'b101011110?01?000?  :  Dest[0] = 1'b1;
	    17'b101011101?00?011?  :  Dest[0] = 1'b1;
	    17'b10101111?0010000?  :  Dest[0] = 1'b1;
	    17'b1010111?000?0111?  :  Dest[0] = 1'b1;
	    17'b?010111?11?00000?  :  Dest[0] = 1'b1;
	    17'b1010111?011??100?  :  Dest[0] = 1'b1;
	    17'b101011101?01?111?  :  Dest[0] = 1'b1;
	    17'b101011110??0111??  :  Dest[0] = 1'b1;
	    17'b1010111011?011?0?  :  Dest[0] = 1'b1;
	    17'b10101111000?1?1??  :  Dest[0] = 1'b1;
	    17'b1010111?0?0110?1?  :  Dest[0] = 1'b1;
	    17'b1010111?100010???  :  Dest[0] = 1'b1;
	    17'b101011110?01?111?  :  Dest[0] = 1'b1;
	    17'b101011101?10?1?1?  :  Dest[0] = 1'b1;
	    17'b?010111010?1??00?  :  Dest[0] = 1'b1;
	    17'b101011111011???0?  :  Dest[0] = 1'b1;
	    17'b00?0?1111????????  :  Dest[0] = 1'b1;
	    17'b10101111000???11?  :  Dest[0] = 1'b1;
	    17'b101011101110?00??  :  Dest[0] = 1'b1;
	    17'b101011110?011??1?  :  Dest[0] = 1'b1;
	    17'b101011100?11000??  :  Dest[0] = 1'b1;
	    17'b1010111?0??01010?  :  Dest[0] = 1'b1;
	    17'b1010111001000????  :  Dest[0] = 1'b1;
	    17'b1010111001?1001??  :  Dest[0] = 1'b1;
	    17'b101011101101?00??  :  Dest[0] = 1'b1;
	    17'b1010111010?1101??  :  Dest[0] = 1'b1;
	    17'b00?0?11000???????  :  Dest[0] = 1'b1;
	    17'b1010111?101?01???  :  Dest[0] = 1'b1;
	    17'b10101111?0001?1??  :  Dest[0] = 1'b1;
	    17'b1010111?01110??0?  :  Dest[0] = 1'b1;
	    17'b1010111?00?001?1?  :  Dest[0] = 1'b1;
	    17'b10101110??0?1001?  :  Dest[0] = 1'b1;
	    17'b1010111011?01?1??  :  Dest[0] = 1'b1;
	    17'b1010111?10110????  :  Dest[0] = 1'b1;
	    17'b1010111?01?11?00?  :  Dest[0] = 1'b1;
	    17'b10101110?00??010?  :  Dest[0] = 1'b1;
	    17'b101011101?0111???  :  Dest[0] = 1'b1;
	    17'b1010111?00?011?0?  :  Dest[0] = 1'b1;
	    17'b1010111?01?0100??  :  Dest[0] = 1'b1;
	    17'b1010111010000????  :  Dest[0] = 1'b1;
	    17'b1010111?00011?0??  :  Dest[0] = 1'b1;
	    17'b1010111?0001?0???  :  Dest[0] = 1'b1;
	    17'b1010111?101??1?1?  :  Dest[0] = 1'b1;
	    17'b1010111?011?11???  :  Dest[0] = 1'b1;
	    17'b1010111?0?101????  :  Dest[0] = 1'b1;
	    17'b1010111??0?010?1?  :  Dest[0] = 1'b1;
	    17'b00001111?1???????  :  Dest[0] = 1'b1;
	    17'b1010111?0?000??0?  :  Dest[0] = 1'b1;
	    17'b1010111?0010?0???  :  Dest[0] = 1'b1;
	    17'b?010011???11?00?0  :  Dest[0] = 1'b1;
	    17'b?110011??1???????  :  Dest[0] = 1'b1;
	    17'b?110011?1????????  :  Dest[0] = 1'b1;
	    17'b?010111111?1?????  :  Dest[0] = 1'b1;
	    17'b0?01111??????????  :  Dest[0] = 1'b1;
	    17'b0?10?11??????????  :  Dest[0] = 1'b1;
	    17'b00?0011??????????  :  Dest[0] = 1'b1;
	    17'b?0101111110??????  :  Dest[0] = 1'b1;
	    17'b110?111??????????  :  Dest[0] = 1'b1;
	    default : Dest[0] = 1'b0;
	endcase
end
endmodule

module autogen_Zb_instr (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcB,
output reg [4:0] Zb_instr
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0]})
	    17'b01100110010000010  :  Zb_instr[4] = 1'b1;
	    17'b001001100101??101  :  Zb_instr[4] = 1'b1;
	    17'b011001100100001?0  :  Zb_instr[4] = 1'b1;
	    17'b00100110110???101  :  Zb_instr[4] = 1'b1;
	    default : Zb_instr[4] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1]})
	    21'b0?1001101100000010010  :  Zb_instr[3] = 1'b1;
	    21'b01100110000100100????  :  Zb_instr[3] = 1'b1;
	    21'b011001101000001?0????  :  Zb_instr[3] = 1'b1;
	    21'b01100110100000111????  :  Zb_instr[3] = 1'b1;
	    21'b01100110110000?01????  :  Zb_instr[3] = 1'b1;
	    default : Zb_instr[3] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0]})
	    17'b011001100001011??  :  Zb_instr[2] = 1'b1;
	    17'b011001101000001?0  :  Zb_instr[2] = 1'b1;
	    17'b011001100100001?0  :  Zb_instr[2] = 1'b1;
	    17'b01100110110000?01  :  Zb_instr[2] = 1'b1;
	    default : Zb_instr[2] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    22'b0?10011011000000100010  :  Zb_instr[1] = 1'b1;
	    22'b0?10011011000000100001  :  Zb_instr[1] = 1'b1;
	    22'b0110011000010111??????  :  Zb_instr[1] = 1'b1;
	    22'b01100110010000010?????  :  Zb_instr[1] = 1'b1;
	    22'b01100110000100100?????  :  Zb_instr[1] = 1'b1;
	    22'b001001100101??101?????  :  Zb_instr[1] = 1'b1;
	    22'b01100110100000111?????  :  Zb_instr[1] = 1'b1;
	    22'b01100110110000?01?????  :  Zb_instr[1] = 1'b1;
	    default : Zb_instr[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    22'b0010011011000000100101  :  Zb_instr[0] = 1'b1;
	    22'b00100110110000001000?0  :  Zb_instr[0] = 1'b1;
	    22'b011001100001011?1?????  :  Zb_instr[0] = 1'b1;
	    22'b01100110100000100?????  :  Zb_instr[0] = 1'b1;
	    22'b01100110010000?10?????  :  Zb_instr[0] = 1'b1;
	    22'b001001101101??101?????  :  Zb_instr[0] = 1'b1;
	    22'b01100110100000111?????  :  Zb_instr[0] = 1'b1;
	    22'b01100110110000101?????  :  Zb_instr[0] = 1'b1;
	    default : Zb_instr[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_rf_rd_op_valid (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] fp_rf_rd_op_valid
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[0]})
	    13'b10?0011?10000  :  fp_rf_rd_op_valid[0] = 1'b1;
	    13'b10?00111?1000  :  fp_rf_rd_op_valid[0] = 1'b1;
	    13'b10?0011000?00  :  fp_rf_rd_op_valid[0] = 1'b1;
	    13'b10?001100?0?0  :  fp_rf_rd_op_valid[0] = 1'b1;
	    13'b0100111??????  :  fp_rf_rd_op_valid[0] = 1'b1;
	    13'b100??11??????  :  fp_rf_rd_op_valid[0] = 1'b1;
	    default : fp_rf_rd_op_valid[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_mad_type_inst (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] fp_mad_type_inst
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[0]})
	    13'b10?0011000?00  :  fp_mad_type_inst[0] = 1'b1;
	    13'b10?00110000?0  :  fp_mad_type_inst[0] = 1'b1;
	    13'b100??11??????  :  fp_mad_type_inst[0] = 1'b1;
	    default : fp_mad_type_inst[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_rf_store_rd_en (
input [6:0] Opcode,
input [2:0] funct3,
output reg [0:0] fp_rf_store_rd_en
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0]})
	    10'b0100111010  :  fp_rf_store_rd_en[0] = 1'b1;
	    10'b0100111001  :  fp_rf_store_rd_en[0] = 1'b1;
	    default : fp_rf_store_rd_en[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_op_int_rs1 (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] fp_op_int_rs1
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[3], funct7[2], funct7[0]})
	    12'b101001111100  :  fp_op_int_rs1[0] = 1'b1;
	    default : fp_op_int_rs1[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_rf_rd_p2_is_rs2 (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] fp_rf_rd_p2_is_rs2
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[0]})
	    12'b101001100000  :  fp_rf_rd_p2_is_rs2[0] = 1'b1;
	    default : fp_rf_rd_p2_is_rs2[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_rd_zero_p2 (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] fp_rd_zero_p2
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[0]})
	    13'b1010011001000  :  fp_rd_zero_p2[0] = 1'b1;
	    13'b1010011000100  :  fp_rd_zero_p2[0] = 1'b1;
	    13'b101001111?000  :  fp_rd_zero_p2[0] = 1'b1;
	    13'b1010011110?00  :  fp_rd_zero_p2[0] = 1'b1;
	    13'b0?00111??????  :  fp_rd_zero_p2[0] = 1'b1;
	    13'b1010011?10000  :  fp_rd_zero_p2[0] = 1'b1;
	    default : fp_rd_zero_p2[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_rd_one_p1 (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] fp_rd_one_p1
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[0]})
	    13'b1010011?10000  :  fp_rd_one_p1[0] = 1'b1;
	    13'b10100110000?0  :  fp_rd_one_p1[0] = 1'b1;
	    13'b101001111?000  :  fp_rd_one_p1[0] = 1'b1;
	    13'b1010011110?00  :  fp_rd_one_p1[0] = 1'b1;
	    13'b0?00111??????  :  fp_rd_one_p1[0] = 1'b1;
	    default : fp_rd_one_p1[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_rd_neg_p1 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] fp_rd_neg_p1
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[0], funct3[2], funct3[1], funct3[0]})
	    16'b1010011001000001  :  fp_rd_neg_p1[0] = 1'b1;
	    16'b1001?11?????????  :  fp_rd_neg_p1[0] = 1'b1;
	    default : fp_rd_neg_p1[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_rd_neg_p2 (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] fp_rd_neg_p2
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[3], funct7[2], funct7[0]})
	    12'b101001100010  :  fp_rd_neg_p2[0] = 1'b1;
	    12'b100?111?????  :  fp_rd_neg_p2[0] = 1'b1;
	    default : fp_rd_neg_p2[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_is_f16 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcB,
output reg [0:0] fp_is_f16
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    22'b10?00111?1001000?00000  :  fp_is_f16[0] = 1'b1;
	    22'b10?0011?100010???00000  :  fp_is_f16[0] = 1'b1;
	    22'b10?001111??01000000000  :  fp_is_f16[0] = 1'b1;
	    22'b10100110100000???00010  :  fp_is_f16[0] = 1'b1;
	    22'b10?0011110?010???0000?  :  fp_is_f16[0] = 1'b1;
	    22'b10?001100?0?1000??????  :  fp_is_f16[0] = 1'b1;
	    22'b10?0011?0100100?0?????  :  fp_is_f16[0] = 1'b1;
	    22'b0?00111???????001?????  :  fp_is_f16[0] = 1'b1;
	    22'b10?0011?01001000??????  :  fp_is_f16[0] = 1'b1;
	    22'b10?00110000?10????????  :  fp_is_f16[0] = 1'b1;
	    22'b10?0011000?010????????  :  fp_is_f16[0] = 1'b1;
	    22'b100??11?????10????????  :  fp_is_f16[0] = 1'b1;
	    default : fp_is_f16[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_take_f16_src (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcB,
output reg [0:0] fp_take_f16_src
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct7[0], funct3[2], funct3[1], funct3[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    22'b10?00111?1001000100000  :  fp_take_f16_src[0] = 1'b1;
	    22'b10100110100000???00010  :  fp_take_f16_src[0] = 1'b1;
	    22'b10?00111100010???0000?  :  fp_take_f16_src[0] = 1'b1;
	    22'b10?001100?0?1000??????  :  fp_take_f16_src[0] = 1'b1;
	    22'b10?0011?0100100?0?????  :  fp_take_f16_src[0] = 1'b1;
	    22'b10?0011?01001000??????  :  fp_take_f16_src[0] = 1'b1;
	    22'b10?0011000?010????????  :  fp_take_f16_src[0] = 1'b1;
	    22'b10?00110000?10????????  :  fp_take_f16_src[0] = 1'b1;
	    22'b100??11?????10????????  :  fp_take_f16_src[0] = 1'b1;
	    default : fp_take_f16_src[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_load_vld (
input [6:0] Opcode,
input [2:0] funct3,
output reg [0:0] fp_load_vld
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0]})
	    10'b0000111010  :  fp_load_vld[0] = 1'b1;
	    10'b0000111001  :  fp_load_vld[0] = 1'b1;
	    default : fp_load_vld[0] = 1'b0;
	endcase
end
endmodule

module autogen_int_to_fp_mov (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] int_to_fp_mov
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[0]})
	    13'b1010011111100  :  int_to_fp_mov[0] = 1'b1;
	    default : int_to_fp_mov[0] = 1'b0;
	endcase
end
endmodule

module autogen_fp_to_int_mov (
input [6:0] Opcode,
input [2:0] funct3,
output reg [0:0] fp_to_int_mov
);

always_comb begin
fp_to_int_mov[0] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for fp_to_int_mov[0]

end
endmodule

module autogen_int_to_fp_cvt (
input [6:0] Opcode,
input [6:0] funct7,
output reg [0:0] int_to_fp_cvt
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[0]})
	    13'b1010011110100  :  int_to_fp_cvt[0] = 1'b1;
	    default : int_to_fp_cvt[0] = 1'b0;
	endcase
end
endmodule

module autogen_out_from_vec_int (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] out_from_vec_int
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111?0?01?100  :  out_from_vec_int[0] = 1'b1;
	    16'b10101110?000001?  :  out_from_vec_int[0] = 1'b1;
	    16'b10101110?0111?00  :  out_from_vec_int[0] = 1'b1;
	    16'b101011111??11?10  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?10000?10  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?010?101?  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?011?0011  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?1000?000  :  out_from_vec_int[0] = 1'b1;
	    16'b101011110?00?011  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111011???100  :  out_from_vec_int[0] = 1'b1;
	    16'b101011111???0110  :  out_from_vec_int[0] = 1'b1;
	    16'b101011110???1?00  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?1101?010  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?01?1?011  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?001?1?00  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111000??0?00  :  out_from_vec_int[0] = 1'b1;
	    16'b10101111??1?1?10  :  out_from_vec_int[0] = 1'b1;
	    16'b10101110??0100?0  :  out_from_vec_int[0] = 1'b1;
	    16'b10101110111??01?  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?011?0?00  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?1??00010  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111011?0?0?0  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111000???010  :  out_from_vec_int[0] = 1'b1;
	    16'b101011110?0???00  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111?010?1??0  :  out_from_vec_int[0] = 1'b1;
	    16'b101011101000010?  :  out_from_vec_int[0] = 1'b1;
	    16'b101011101011110?  :  out_from_vec_int[0] = 1'b1;
	    16'b101011100111?10?  :  out_from_vec_int[0] = 1'b1;
	    16'b101011101?00?011  :  out_from_vec_int[0] = 1'b1;
	    16'b101011101?11101?  :  out_from_vec_int[0] = 1'b1;
	    16'b101011110?1?101?  :  out_from_vec_int[0] = 1'b1;
	    16'b101011100?01101?  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111110????10  :  out_from_vec_int[0] = 1'b1;
	    16'b101011101?0???00  :  out_from_vec_int[0] = 1'b1;
	    16'b10101111?01???10  :  out_from_vec_int[0] = 1'b1;
	    16'b1010111001?1?1?0  :  out_from_vec_int[0] = 1'b1;
	    16'b10101110010???10  :  out_from_vec_int[0] = 1'b1;
	    default : out_from_vec_int[0] = 1'b0;
	endcase
end
endmodule

module autogen_vfp_mad_type_inst (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] vfp_mad_type_inst
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b10101111?1?00?01  :  vfp_mad_type_inst[0] = 1'b1;
	    16'b10101110000?0?01  :  vfp_mad_type_inst[0] = 1'b1;
	    16'b101011110?111101  :  vfp_mad_type_inst[0] = 1'b1;
	    16'b1010111110??0?01  :  vfp_mad_type_inst[0] = 1'b1;
	    16'b1010111101????01  :  vfp_mad_type_inst[0] = 1'b1;
	    16'b10101111?11???01  :  vfp_mad_type_inst[0] = 1'b1;
	    16'b10101111??100?01  :  vfp_mad_type_inst[0] = 1'b1;
	    default : vfp_mad_type_inst[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_wdeop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
output reg [0:0] v_wdeop
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], SrcA[4], SrcA[3], SrcA[2], SrcA[1], SrcA[0]})
	    21'b101011111??00?10?????  :  v_wdeop[0] = 1'b1;
	    21'b101011111?1?1?10?????  :  v_wdeop[0] = 1'b1;
	    21'b101011111?01??10?????  :  v_wdeop[0] = 1'b1;
	    21'b101011111???0110?????  :  v_wdeop[0] = 1'b1;
	    21'b1010111?1001000101??0  :  v_wdeop[0] = 1'b1;
	    21'b1010111?10010001010??  :  v_wdeop[0] = 1'b1;
	    21'b1010111?1001000101?1?  :  v_wdeop[0] = 1'b1;
	    21'b10101111111???01?????  :  v_wdeop[0] = 1'b1;
	    21'b1010111110????10?????  :  v_wdeop[0] = 1'b1;
	    21'b101011111??00?01?????  :  v_wdeop[0] = 1'b1;
	    21'b1010111110??0?01?????  :  v_wdeop[0] = 1'b1;
	    default : v_wdeop[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_nrwop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
output reg [0:0] v_nrwop
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], SrcA[4], SrcA[3]})
	    18'b101011101001000110  :  v_nrwop[0] = 1'b1;
	    18'b10101111011???00??  :  v_nrwop[0] = 1'b1;
	    18'b10101111011??011??  :  v_nrwop[0] = 1'b1;
	    default : v_nrwop[0] = 1'b0;
	endcase
end
endmodule

module autogen_vfp_rf_rd_op_valid (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
input [4:0] SrcB,
output reg [0:0] vfp_rf_rd_op_valid
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], SrcA[4], SrcA[3], SrcA[2], SrcA[1], SrcA[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b1010111?1?000101?????00000  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?1001?00110000?????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?1001000101??0?????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b10101110??00000100000?????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?100100010?0???????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?100100010??1??????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?1001000110????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?1110?101??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111??1111101??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?0100??01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b101011100??10101??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?00100?01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b101011100?0?0?01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b101011101?111101?????00000  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b10101111?11???01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b101011110?111101??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111101????01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111000???001??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111110??0?01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b10101111100??001??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b10101110110?1?01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    26'b1010111?11?00?01??????????  :  vfp_rf_rd_op_valid[0] = 1'b1;
	    default : vfp_rf_rd_op_valid[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_src1hw (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_src1hw
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[1], funct3[1], funct3[0]})
	    14'b10101111101001  :  v_src1hw[0] = 1'b1;
	    14'b10101111101?10  :  v_src1hw[0] = 1'b1;
	    default : v_src1hw[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_rf_store_rd_en (
input [6:0] Opcode,
input [2:0] funct3,
output reg [0:0] v_rf_store_rd_en
);

always_comb begin
v_rf_store_rd_en[0] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_rf_store_rd_en[0]

end
endmodule

module autogen_v_math_fmt (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [3:0] v_math_fmt
);

always_comb begin
v_math_fmt[3] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_math_fmt[3]

v_math_fmt[2] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_math_fmt[2]

v_math_fmt[1] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_math_fmt[1]

v_math_fmt[0] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_math_fmt[0]

end
endmodule

module autogen_v_rf_rd_p2_is_rs2 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_rf_rd_p2_is_rs2
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b10101111010?1?10  :  v_rf_rd_p2_is_rs2[0] = 1'b1;
	    16'b1010111000??1001  :  v_rf_rd_p2_is_rs2[0] = 1'b1;
	    16'b1010111110??0?01  :  v_rf_rd_p2_is_rs2[0] = 1'b1;
	    16'b1010111100111101  :  v_rf_rd_p2_is_rs2[0] = 1'b1;
	    16'b10101110000?0?01  :  v_rf_rd_p2_is_rs2[0] = 1'b1;
	    16'b10101111010???01  :  v_rf_rd_p2_is_rs2[0] = 1'b1;
	    16'b10101111100??001  :  v_rf_rd_p2_is_rs2[0] = 1'b1;
	    default : v_rf_rd_p2_is_rs2[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_acc_val (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_acc_val
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b10101110000?0?01  :  v_acc_val[0] = 1'b1;
	    16'b10101111111??110  :  v_acc_val[0] = 1'b1;
	    16'b1010111000??1001  :  v_acc_val[0] = 1'b1;
	    16'b1010111101??1?10  :  v_acc_val[0] = 1'b1;
	    16'b101011111110??10  :  v_acc_val[0] = 1'b1;
	    16'b10101111?11?1?10  :  v_acc_val[0] = 1'b1;
	    16'b1010111110??0?01  :  v_acc_val[0] = 1'b1;
	    16'b10101111100??001  :  v_acc_val[0] = 1'b1;
	    16'b101011110?111101  :  v_acc_val[0] = 1'b1;
	    16'b1010111101????01  :  v_acc_val[0] = 1'b1;
	    16'b10101111?11???01  :  v_acc_val[0] = 1'b1;
	    default : v_acc_val[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_rd_onep1 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_rd_onep1
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111100111101  :  v_rd_onep1[0] = 1'b1;
	    16'b10101110000??001  :  v_rd_onep1[0] = 1'b1;
	    16'b10101110000?0?01  :  v_rd_onep1[0] = 1'b1;
	    16'b1010111110??0?01  :  v_rd_onep1[0] = 1'b1;
	    16'b10101111100??001  :  v_rd_onep1[0] = 1'b1;
	    default : v_rd_onep1[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_rd_zerop2 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_rd_zerop2
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[1], funct3[0]})
	    15'b101011111100001  :  v_rd_zerop2[0] = 1'b1;
	    15'b101011110010001  :  v_rd_zerop2[0] = 1'b1;
	    default : v_rd_zerop2[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_rf_rdneg0 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_rf_rdneg0
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[1], funct3[0]})
	    15'b101011100001001  :  v_rf_rdneg0[0] = 1'b1;
	    15'b1010111110?1001  :  v_rf_rdneg0[0] = 1'b1;
	    15'b1010111101??101  :  v_rf_rdneg0[0] = 1'b1;
	    15'b10101111?11?101  :  v_rf_rdneg0[0] = 1'b1;
	    default : v_rf_rdneg0[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_rd_neg1 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_rd_neg1
);

always_comb begin
v_rd_neg1[0] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_rd_neg1[0]

end
endmodule

module autogen_v_rd_neg2 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_rd_neg2
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111100111101  :  v_rd_neg2[0] = 1'b1;
	    16'b1010111101?10?01  :  v_rd_neg2[0] = 1'b1;
	    16'b10101111?1110?01  :  v_rd_neg2[0] = 1'b1;
	    16'b1010111101?01?01  :  v_rd_neg2[0] = 1'b1;
	    16'b10101111?1101?01  :  v_rd_neg2[0] = 1'b1;
	    default : v_rd_neg2[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_cmpmul (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_cmpmul
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[2], funct7[1], funct3[1], funct3[0]})
	    14'b10101111011110  :  v_cmpmul[0] = 1'b1;
	    default : v_cmpmul[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_rnden (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_rnden
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b101011110?111?00  :  v_rnden[0] = 1'b1;
	    16'b10101110010???10  :  v_rnden[0] = 1'b1;
	    16'b1010111101?1?011  :  v_rnden[0] = 1'b1;
	    16'b1010111101?1??00  :  v_rnden[0] = 1'b1;
	    default : v_rnden[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_saturate (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_saturate
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct3[2], funct3[1], funct3[0]})
	    15'b101011110000011  :  v_saturate[0] = 1'b1;
	    15'b10101111000??00  :  v_saturate[0] = 1'b1;
	    default : v_saturate[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_mulh (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_mulh
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[1], funct3[0]})
	    15'b10101111001?010  :  v_mulh[0] = 1'b1;
	    15'b101011110011?10  :  v_mulh[0] = 1'b1;
	    default : v_mulh[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_usemask (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [0:0] vm,
output reg [0:0] v_usemask
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct3[2], funct3[1], funct3[0], vm[0]})
	    16'b1010111010000110  :  v_usemask[0] = 1'b1;
	    16'b10101110100??000  :  v_usemask[0] = 1'b1;
	    default : v_usemask[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_wrmask (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_wrmask
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111010001011  :  v_wrmask[0] = 1'b1;
	    16'b10101110100?1?00  :  v_wrmask[0] = 1'b1;
	    default : v_wrmask[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_inversesub (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_inversesub
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111000011100  :  v_inversesub[0] = 1'b1;
	    16'b1010111000011011  :  v_inversesub[0] = 1'b1;
	    default : v_inversesub[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_issgn_src2 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_issgn_src2
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b10101111?0001000  :  v_issgn_src2[0] = 1'b1;
	    16'b1010111000000010  :  v_issgn_src2[0] = 1'b1;
	    16'b1010111111?10110  :  v_issgn_src2[0] = 1'b1;
	    16'b10101110010?1?10  :  v_issgn_src2[0] = 1'b1;
	    16'b101011111101??10  :  v_issgn_src2[0] = 1'b1;
	    16'b1010111100001011  :  v_issgn_src2[0] = 1'b1;
	    16'b1010111101?11011  :  v_issgn_src2[0] = 1'b1;
	    16'b1010111?001?1010  :  v_issgn_src2[0] = 1'b1;
	    16'b101011110011??10  :  v_issgn_src2[0] = 1'b1;
	    16'b10101111000?1?00  :  v_issgn_src2[0] = 1'b1;
	    16'b101011110??11?00  :  v_issgn_src2[0] = 1'b1;
	    16'b101011111?101?10  :  v_issgn_src2[0] = 1'b1;
	    16'b1010111110??1?10  :  v_issgn_src2[0] = 1'b1;
	    16'b10101111?01?1?10  :  v_issgn_src2[0] = 1'b1;
	    default : v_issgn_src2[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_issgn_src1 (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_issgn_src1
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b10101111?0001000  :  v_issgn_src1[0] = 1'b1;
	    16'b1010111100?11?00  :  v_issgn_src1[0] = 1'b1;
	    16'b1010111000000010  :  v_issgn_src1[0] = 1'b1;
	    16'b10101110010?1?10  :  v_issgn_src1[0] = 1'b1;
	    16'b1010111101011011  :  v_issgn_src1[0] = 1'b1;
	    16'b1010111100001011  :  v_issgn_src1[0] = 1'b1;
	    16'b101011110?011?00  :  v_issgn_src1[0] = 1'b1;
	    16'b1010111?001?1010  :  v_issgn_src1[0] = 1'b1;
	    16'b101011111?1?1?10  :  v_issgn_src1[0] = 1'b1;
	    16'b10101111000?1?00  :  v_issgn_src1[0] = 1'b1;
	    16'b101011111??11?10  :  v_issgn_src1[0] = 1'b1;
	    16'b1010111110??1?10  :  v_issgn_src1[0] = 1'b1;
	    16'b10101111?01?1?10  :  v_issgn_src1[0] = 1'b1;
	    default : v_issgn_src1[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_cryorbrw (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_cryorbrw
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct3[2], funct3[1], funct3[0]})
	    15'b101011101000011  :  v_cryorbrw[0] = 1'b1;
	    15'b10101110100??00  :  v_cryorbrw[0] = 1'b1;
	    default : v_cryorbrw[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_addorsub (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_addorsub
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111?00010?00  :  v_addorsub[0] = 1'b1;
	    16'b1010111?0001?100  :  v_addorsub[0] = 1'b1;
	    16'b10101110001??010  :  v_addorsub[0] = 1'b1;
	    16'b1010111000011011  :  v_addorsub[0] = 1'b1;
	    16'b101011100101??10  :  v_addorsub[0] = 1'b1;
	    16'b1010111110?1??10  :  v_addorsub[0] = 1'b1;
	    16'b101011110001??00  :  v_addorsub[0] = 1'b1;
	    16'b101011101001??00  :  v_addorsub[0] = 1'b1;
	    default : v_addorsub[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_avg (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_avg
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct3[1], funct3[0]})
	    13'b1010111001010  :  v_avg[0] = 1'b1;
	    default : v_avg[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_imulop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_imulop
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b10101111110?0?10  :  v_imulop[0] = 1'b1;
	    16'b10101111?1?11?10  :  v_imulop[0] = 1'b1;
	    16'b101011111110??10  :  v_imulop[0] = 1'b1;
	    16'b1010111111??0110  :  v_imulop[0] = 1'b1;
	    16'b1010111100111??0  :  v_imulop[0] = 1'b1;
	    16'b10101111001???10  :  v_imulop[0] = 1'b1;
	    16'b1010111101??1?10  :  v_imulop[0] = 1'b1;
	    default : v_imulop[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_iaddop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_iaddop
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111?0001?100  :  v_iaddop[0] = 1'b1;
	    16'b1010111?1000?000  :  v_iaddop[0] = 1'b1;
	    16'b101011100000001?  :  v_iaddop[0] = 1'b1;
	    16'b1010111?000?0?00  :  v_iaddop[0] = 1'b1;
	    16'b10101110010???10  :  v_iaddop[0] = 1'b1;
	    16'b1010111110????10  :  v_iaddop[0] = 1'b1;
	    16'b1010111000011011  :  v_iaddop[0] = 1'b1;
	    16'b101011110000?011  :  v_iaddop[0] = 1'b1;
	    16'b101011101000?011  :  v_iaddop[0] = 1'b1;
	    16'b10101110001??010  :  v_iaddop[0] = 1'b1;
	    16'b10101111000???00  :  v_iaddop[0] = 1'b1;
	    16'b10101110100???00  :  v_iaddop[0] = 1'b1;
	    default : v_iaddop[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_fp_sel_scalar (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_fp_sel_scalar
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111??1111101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b1010111?0100?101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b1010111?00100101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b10101111?11??101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b10101110??000101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b1010111?11?00101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b101011100??10101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b101011101?111101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b101011110?111101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b1010111110??0101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b1010111011??1101  :  v_fp_sel_scalar[0] = 1'b1;
	    16'b1010111101???101  :  v_fp_sel_scalar[0] = 1'b1;
	    default : v_fp_sel_scalar[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_sel_scalar (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [0:0] vm,
output reg [0:0] v_sel_scalar
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], vm[0]})
	    17'b101011101?0??1000  :  v_sel_scalar[0] = 1'b1;
	    17'b10101111??1?1110?  :  v_sel_scalar[0] = 1'b1;
	    17'b10101111?1?11110?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111000??0100?  :  v_sel_scalar[0] = 1'b1;
	    17'b101011110???1100?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111?010?11?0?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111?011?0100?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111?001?1100?  :  v_sel_scalar[0] = 1'b1;
	    17'b101011110?0??100?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111010000101?  :  v_sel_scalar[0] = 1'b1;
	    17'b10101110???11100?  :  v_sel_scalar[0] = 1'b1;
	    17'b101011100111?10??  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111110???110?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111?10000110?  :  v_sel_scalar[0] = 1'b1;
	    17'b101011111???0110?  :  v_sel_scalar[0] = 1'b1;
	    17'b10101111?01??110?  :  v_sel_scalar[0] = 1'b1;
	    17'b10101110010??110?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111011???100?  :  v_sel_scalar[0] = 1'b1;
	    17'b101011101?0?1100?  :  v_sel_scalar[0] = 1'b1;
	    17'b1010111001?1?1?0?  :  v_sel_scalar[0] = 1'b1;
	    default : v_sel_scalar[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_sel_imm (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_sel_imm
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111011?0?011  :  v_sel_imm[0] = 1'b1;
	    16'b1010111?00000011  :  v_sel_imm[0] = 1'b1;
	    16'b1010111?010?1011  :  v_sel_imm[0] = 1'b1;
	    16'b1010111101???011  :  v_sel_imm[0] = 1'b1;
	    16'b10101110?11?0011  :  v_sel_imm[0] = 1'b1;
	    16'b101011101?111011  :  v_sel_imm[0] = 1'b1;
	    16'b101011101?00?011  :  v_sel_imm[0] = 1'b1;
	    16'b101011110??01011  :  v_sel_imm[0] = 1'b1;
	    16'b101011100?011011  :  v_sel_imm[0] = 1'b1;
	    16'b1010111?01?1?011  :  v_sel_imm[0] = 1'b1;
	    default : v_sel_imm[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_shftop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_shftop
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b101011110?101011  :  v_shftop[0] = 1'b1;
	    16'b101011110?101?00  :  v_shftop[0] = 1'b1;
	    16'b1010111101???011  :  v_shftop[0] = 1'b1;
	    16'b1010111101????00  :  v_shftop[0] = 1'b1;
	    default : v_shftop[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_permuteop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_permuteop
);

always_comb begin
v_permuteop[0] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_permuteop[0]

end
endmodule

module autogen_v_p1_dest (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_p1_dest
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct3[1], funct3[0]})
	    13'b1010111101001  :  v_p1_dest[0] = 1'b1;
	    default : v_p1_dest[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_sat_instrn (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_sat_instrn
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct3[2], funct3[1], funct3[0]})
	    15'b101011110000011  :  v_sat_instrn[0] = 1'b1;
	    15'b10101111000??00  :  v_sat_instrn[0] = 1'b1;
	    default : v_sat_instrn[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_bitwiseop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [0:0] vm,
input [4:0] SrcB,
output reg [0:0] v_bitwiseop
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], vm[0]})
	    17'b10101110?1001011?  :  v_bitwiseop[0] = 1'b1;
	    17'b1010111011???010?  :  v_bitwiseop[0] = 1'b1;
	    17'b1010111011?0??00?  :  v_bitwiseop[0] = 1'b1;
	    17'b101011101?1110110  :  v_bitwiseop[0] = 1'b1;
	    17'b10101110?0111?000  :  v_bitwiseop[0] = 1'b1;
	    17'b1010111010111101?  :  v_bitwiseop[0] = 1'b1;
	    17'b10101110001???00?  :  v_bitwiseop[0] = 1'b1;
	    17'b101011100101?011?  :  v_bitwiseop[0] = 1'b1;
	    17'b101011100001?010?  :  v_bitwiseop[0] = 1'b1;
	    17'b1010111011?0?01??  :  v_bitwiseop[0] = 1'b1;
	    17'b10101110000?1010?  :  v_bitwiseop[0] = 1'b1;
	    17'b10101110111??01??  :  v_bitwiseop[0] = 1'b1;
	    17'b10101110?101??00?  :  v_bitwiseop[0] = 1'b1;
	    17'b10101110?10?1?00?  :  v_bitwiseop[0] = 1'b1;
	    17'b1010111011???100?  :  v_bitwiseop[0] = 1'b1;
	    default : v_bitwiseop[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_iterate (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
output reg [0:0] v_iterate
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b10101111100?1001  :  v_iterate[0] = 1'b1;
	    16'b101011111000?000  :  v_iterate[0] = 1'b1;
	    16'b101011100111?10?  :  v_iterate[0] = 1'b1;
	    16'b10101110011?0?00  :  v_iterate[0] = 1'b1;
	    16'b10101110?0010010  :  v_iterate[0] = 1'b1;
	    16'b101011100111?1?0  :  v_iterate[0] = 1'b1;
	    16'b1010111000??1001  :  v_iterate[0] = 1'b1;
	    16'b10101110011?0011  :  v_iterate[0] = 1'b1;
	    16'b10101110?0111010  :  v_iterate[0] = 1'b1;
	    16'b1010111000???010  :  v_iterate[0] = 1'b1;
	    16'b101011100111?011  :  v_iterate[0] = 1'b1;
	    default : v_iterate[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_reductop (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
output reg [0:0] v_reductop
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b101011111000?000  :  v_reductop[0] = 1'b1;
	    16'b10101111100?1001  :  v_reductop[0] = 1'b1;
	    16'b1010111000???010  :  v_reductop[0] = 1'b1;
	    16'b1010111000??1001  :  v_reductop[0] = 1'b1;
	    default : v_reductop[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_onecycle_iterate (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
output reg [0:0] v_onecycle_iterate
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b101011111000?000  :  v_onecycle_iterate[0] = 1'b1;
	    16'b10101111100?1001  :  v_onecycle_iterate[0] = 1'b1;
	    16'b10101110?0010010  :  v_onecycle_iterate[0] = 1'b1;
	    16'b1010111000??1001  :  v_onecycle_iterate[0] = 1'b1;
	    16'b1010111000???010  :  v_onecycle_iterate[0] = 1'b1;
	    16'b10101110?0111010  :  v_onecycle_iterate[0] = 1'b1;
	    default : v_onecycle_iterate[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_vmvgrp (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
output reg [0:0] v_vmvgrp
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], SrcA[4], SrcA[3], SrcA[2], SrcA[1], SrcA[0]})
	    21'b10101111001110110000?  :  v_vmvgrp[0] = 1'b1;
	    21'b101011110011101100?11  :  v_vmvgrp[0] = 1'b1;
	    default : v_vmvgrp[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_scalar_dest (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
output reg [0:0] v_scalar_dest
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0]})
	    16'b1010111010000010  :  v_scalar_dest[0] = 1'b1;
	    16'b1010111010000001  :  v_scalar_dest[0] = 1'b1;
	    default : v_scalar_dest[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_mask_only (
input [6:0] Opcode,
input [6:0] funct7,
input [2:0] funct3,
input [4:0] SrcA,
output reg [0:0] v_mask_only
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct7[6], funct7[5], funct7[4], funct7[3], funct7[2], funct7[1], funct3[2], funct3[1], funct3[0], SrcA[4], SrcA[3], SrcA[2], SrcA[1], SrcA[0]})
	    21'b1010111011?0?01??????  :  v_mask_only[0] = 1'b1;
	    21'b1010111011?0??00?????  :  v_mask_only[0] = 1'b1;
	    21'b1010111011?00?0??????  :  v_mask_only[0] = 1'b1;
	    21'b10101110110??0?0?????  :  v_mask_only[0] = 1'b1;
	    21'b101011101?1000100001?  :  v_mask_only[0] = 1'b1;
	    21'b101011101?100010000?1  :  v_mask_only[0] = 1'b1;
	    21'b101011101?0?1?00?????  :  v_mask_only[0] = 1'b1;
	    21'b101011101?001011?????  :  v_mask_only[0] = 1'b1;
	    21'b1010111011??110??????  :  v_mask_only[0] = 1'b1;
	    21'b10101110111??01??????  :  v_mask_only[0] = 1'b1;
	    21'b1010111011???100?????  :  v_mask_only[0] = 1'b1;
	    21'b10101110110?1?0??????  :  v_mask_only[0] = 1'b1;
	    default : v_mask_only[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_ldst_iterations (
input [6:0] Opcode,
input [2:0] funct3,
input [2:0] sew,
input [2:0] lmul,
input [1:0] mop,
input [2:0] nf,
input [4:0] SrcB,
output reg [5:0] v_ldst_iterations
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    25'b000011111100?011000010000  :  v_ldst_iterations[5] = 1'b1;
	    25'b0?00111111000000?11??????  :  v_ldst_iterations[5] = 1'b1;
	    default : v_ldst_iterations[5] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    25'b00001111110?0011000010000  :  v_ldst_iterations[4] = 1'b1;
	    25'b000011111100?011000010000  :  v_ldst_iterations[4] = 1'b1;
	    25'b0?00111110000001?101?????  :  v_ldst_iterations[4] = 1'b1;
	    25'b0?00111111001001?101?????  :  v_ldst_iterations[4] = 1'b1;
	    25'b0?00111110000000?11??????  :  v_ldst_iterations[4] = 1'b1;
	    25'b0?00111111001000?11??????  :  v_ldst_iterations[4] = 1'b1;
	    25'b0?00111111000111?11??????  :  v_ldst_iterations[4] = 1'b1;
	    25'b0?00111111000000?1?1?????  :  v_ldst_iterations[4] = 1'b1;
	    default : v_ldst_iterations[4] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    25'b00001111110??011000010000  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111110001010?1001????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111010010?1001????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111101000010?1001????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111110001001?101?????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111010001?101?????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111101000001?101?????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111110000001?10?1????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111001001?10?1????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111110001000?11??????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111110000111?11??????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111001111?11??????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111000110?11??????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111010000?11??????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111101000000?11??????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111110000000?1?1?????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111001000?1?1?????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111000111?1?1?????  :  v_ldst_iterations[3] = 1'b1;
	    25'b0?00111111000000?1??1????  :  v_ldst_iterations[3] = 1'b1;
	    default : v_ldst_iterations[3] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b010011111?0011?100100?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?????0011101000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111000001010?001??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b00001111?10?????0011101000  :  v_ldst_iterations[2] = 1'b1;
	    26'b000011111?0?????0011101000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100000001???001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111101010011??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100000?011??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111000111??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111010001??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111101000001??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100?1010?001??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1010010?001??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?011011??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?010010??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?001001??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111101?010??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110100?010??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?000000??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000110???01???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111110000111??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111100?000??001?0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111001111??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111000110??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000000?1??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?0011??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010110?0?01???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100001?0?0?01???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?100??01???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100001?00??01???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111001100??01???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000010101001??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b000011111?0011?110110?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000001?1??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?0111??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100010?0??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1011011??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1001001??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1000000??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100?0001??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110?1001??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110?0000??01??0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110101?00??01???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111000000011??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100000?11???1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1011000??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100000001?1?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010?1000??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000??000??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010100111?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111001?000??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100000?0111?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110001111?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110100011?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010000011?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100?111???1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100?10101001??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0?1110??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111011011??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111010010??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111101000010??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?101011???1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?10100101001??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0110111?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0101?1??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100??110??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0100101?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111001001??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?101?111??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111000000??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110100?11???1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0010011?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111101?0101?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110100?0101?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0000001?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?100?101??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?00?101??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000110??101???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110??101??1???0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100001111?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111100?0001?001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110011111?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110001101?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000000?11?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?00111?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010110?0101???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100001?0?0101???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?100?101???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100001?00?101???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111001100?101???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111110000001??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111110001010??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111010001?10?1?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111101000001?10?1?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111110010011??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000??01??1001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111101001011??????0000  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?01?010?1001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000001?1?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000001?11?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010??010?1001?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?01111?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100010?01?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?10110111?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111110000111?1?1??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111001111?1?1??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?10010011?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111000110?1?1??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?10000001?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?001001?10?1?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100?00011?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110?10011?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110?00001?01??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110101?00?101???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111000111?1??1?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100000?11??11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000000111?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100011?1?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011100000?11?1?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1011000?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?10110001?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000?0?11?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010?1000?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000??000?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110101?000?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010?10001?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000??0001?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111001?000?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111001?0001?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000??0?1?101??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110101?0?1?101??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111001?0?1?101??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?10?1001?101??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100010?0?1?1??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1000000?1?1??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110?0000?1?1??????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?000000?1??1?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0?1110?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100?111?1?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0?11101?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111010010?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110110111?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111101000010?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?101011??11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110100101?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010000101?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111100?000?1??1?????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?101011?1?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100??110?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111001001?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0101?11?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100??1101?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111111000000?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110010011?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?101?1111?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110000001?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110100?11??11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010??111?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?0?0101?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110100?11?1?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?100?101?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?100?1011?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?00?1011?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110??101?11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111110??1011?1???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111110001010?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100010101?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001110000??011?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100100111?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010010111?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111?01?11??11???????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?00111110000001?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111100000011?????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111?1011011?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?001111010?1011?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011110101?011?1????????  :  v_ldst_iterations[2] = 1'b1;
	    26'b0?0011111001?011?1????????  :  v_ldst_iterations[2] = 1'b1;
	    default : v_ldst_iterations[2] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b00001111110??01100001?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?????00?1101000  :  v_ldst_iterations[1] = 1'b1;
	    26'b00001111?10?????00?1101000  :  v_ldst_iterations[1] = 1'b1;
	    26'b000011111?0?????00?1101000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000000?1??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?0011??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100001?00??0?1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?10?1?0?1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b000011111?0011?110110?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100?1001?0?1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000001?1???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?0111???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?1011011??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?1010010??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000?01???0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?000111??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100011???0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?1001001??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?1000000??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100?0001??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110?1001??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100?111??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110?0000??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110101?00??0?1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100001?0?0???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000?11????1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000??000???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111001?000???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?01?010??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?00?000??0?1?0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000001???????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000?011??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111111000111??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100?111????1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0?1110???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?101011????1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10110?0???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0101?1???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100??110???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?101?111???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111101010011??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110100?11????1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10?1000???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?100?101???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111111010001??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?00?101???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111101000001??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110??101???1??0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000000?11?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?00111?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111110000001??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?010010??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100001?00?10?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111110001010??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?10?110?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111101?010??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?000000??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111110010011??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111101001011??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100?000??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100?100110?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?011011??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000001?1?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000001?11??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?01111??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?001001??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110100?010??????0000  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10110111?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10100101?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000?01?1?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0001111?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0100011?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100011?1?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10010011?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10000001?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110?10011?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100?1111?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110?00001?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110101?00?10?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?1001110?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100001?0?01??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100011?1?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000?11?1??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000?0?11?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000??0001??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111001?0001??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000??0?1?10?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?01?0101?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?01?001?10?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010??001?10?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?000111?1??1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?00?0001?0?1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100011??1??1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?1000000?1??1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000001?1?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100?111?1??1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110?0000?1??1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000?0111?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111111000111?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111111010001?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110001111?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111101000001?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100?111?1??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0?11101??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110100011?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?101011?1??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100??110?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011100000??1??1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10110?01??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0101?11??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010?011??1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100??1101??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000??0?0?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?101?1111??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110101?0?0?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010100111?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111001?0?0?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10?1000?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010??111?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0?0101?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110100?11?1??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?10?10001??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?100?101?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?100?1011??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?00?1011??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010000011?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110??101?1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111110??1011??1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0100101?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?00?000?1??1?????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111110001010?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100010101?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?000000?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111101?0101?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0000001?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100100111?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010010111?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100?000?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?01?11??1?1??????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111100?0001?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?00111110000001?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0110111?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111100000011?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?001001?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?0010011?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110100?0101?????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111?1011011?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010?1011?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011110101?011?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111001?011?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001110000??01??1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?0011111?01?010?1????????  :  v_ldst_iterations[1] = 1'b1;
	    26'b0?001111010??010?1????????  :  v_ldst_iterations[1] = 1'b1;
	    default : v_ldst_iterations[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b00001111110??01100001?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000?????000?101000  :  v_ldst_iterations[0] = 1'b1;
	    26'b00001111?10?????0011101000  :  v_ldst_iterations[0] = 1'b1;
	    26'b000011111?0?????0011101000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000?????00?1101000  :  v_ldst_iterations[0] = 1'b1;
	    26'b00001111?10?????000?101000  :  v_ldst_iterations[0] = 1'b1;
	    26'b000011111?0?????000?101000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111000000??1????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000?0?11????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000000?1??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000?0011??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011100000??1?????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111101010011??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111111010001??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111101000001??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?1011011??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?1010010??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011100000?01???????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?000111??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111100011???????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?1001001??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?1000000??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111100?0001??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110?1001??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111100?111??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111110001010??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110?0000??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111110010011??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111101001011??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?011011??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10?011?????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000??0??????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0?01?1????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?001001??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?100?11?????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011110100?010??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?100?1?1????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10??111????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?101?00?????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?00?1?1????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010??0?0????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110??1?1????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111100??00?????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?01?010??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?00?000??????0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111000000??1?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000?0?11?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111000000??11???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000?0?111???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0??11?????1?0000  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000000?11?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000?00111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011100000??1??1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011100000??1?1???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010100111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010000011?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10110111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10100101?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?000111?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011100000?01?1?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111100011??1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0001111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0100011?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111100011?1?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?1000000?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10010011?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10000001?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111100?111?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111110001010?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110?0000?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110?10011?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111100?1111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111100010101?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110?00001?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111100100111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010010111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?00111110000001?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0110111?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111100000011?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10?011??1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000??0???1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10?011?1???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0?01?1?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?001001?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000??0??1???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0?01?11???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?100?11??1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0010011?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?100?1?1?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10??111?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?100?11?1???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?00?1?1?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011110100?0101?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?100?1?11???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10??1111???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?101?00?1???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?00?1?11???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?01?00?1???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110??1?1?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010??0?01???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111110??1?11???1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000??0?1?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?10??000?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0??000?1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?01?0101?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?01?001?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010??001?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111?1011011?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?00?000?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?00?0001?????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010?1011?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011110101?011?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111001?011?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001110000??01??1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?01?010?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?001111010??010?1????????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0??11??1??1?????  :  v_ldst_iterations[0] = 1'b1;
	    26'b0?0011111?0??11?1???1?????  :  v_ldst_iterations[0] = 1'b1;
	    default : v_ldst_iterations[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_ldst_dest_incr (
input [6:0] Opcode,
input [2:0] funct3,
input [2:0] sew,
input [2:0] lmul,
input [1:0] mop,
input [2:0] nf,
input [4:0] SrcB,
output reg [7:0] v_ldst_dest_incr
);

always_comb begin
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b0?00111000001010?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111000110?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110000111?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111001111?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111010001?0001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111101000001?0001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111000111?0001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001100??0111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010110?0?0111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100010?0?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100001?0?0?0111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?1000000?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?100??0111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000110???0111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100?1010?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100001?00??0111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?1010010?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110?0000?0011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?000000?0001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000001?1??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?0111??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?001001?0001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100?000?0001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000000?1??011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?1011000??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?0011??011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001?000??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111101010011??001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010?1000??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000001???001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100011?1??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110101?00??0111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000?011??001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000??000??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?????0011101000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000101010011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000?11???111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100100?1??011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b000011111?0?????0011101000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?1011011??011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110110?1??011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b00001111?10?????0011101000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010010?1??011?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?011011??001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001001???001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111101101???001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110100101???001?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0?1110??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100??110??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0?0101??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?101011???111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100011010011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?100?101??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?101?111??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110??101??111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111000011110011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110100?11???111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100111110011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111101000110001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110100000110001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100011110001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001100?10111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010110?010111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111000000?0????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100010?010011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100001?0?010111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?100000010011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?100?10111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000110??10111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100?101010011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?01?11???111?0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100001?00?10111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?101001010011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111001001?0????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110?000010011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?00000010001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000001?1?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000001?11?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?01111?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?00100110001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100?00010001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111000000011??????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000000?11?011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?10110001?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?00111?011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001?0001?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010100111?001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010?10001?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000001?1?001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100011??1?11?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111101000010?0????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000??000?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100011?11?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110101?00?10111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000?0111?001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000??0001?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?000111?1?11?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100?111?1?11?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000?0?11?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110001001?101??????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110010011??????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000?11??1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110001001?10?1?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111011011??????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011100000?11?1?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111010001?101??????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100100?11?011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111101001011??????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?10110111?011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110110?11?011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111010001?10?1?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111101000001?101??????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010010?11?011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111101000001?10?1?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0110111?001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001001?1?001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111101101?1?001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0??000?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110100101?1?001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0?11101?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100010?0?1?11?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0?01?1?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110100?0?1?11?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?10?011??1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100??1101?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0?01011?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?10??000?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?00?1?1?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?101011?1?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010000?0?1?11?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?100?1?1?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?100?1011?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110??1?1?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111000111?1?1??????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111000111?1??1?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?101?1111?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110??1011?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?10110?1?1011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?100?11??1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110100?11?1?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?10??111?1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001?0?1?1011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010?10?1?1011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110101?0?1?1011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?101101??1001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000??0?1?1011?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001?01??1001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010?101??1001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111000000?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110101?01??1001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111000110?11???????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100000010????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111000000??1?1??????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000??01??1001?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110000001?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?000111?11???????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100100??1?1??????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111001001?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111000000??1??1?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100100??1??1?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111001111?11???????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?01?11?1?111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111100100110????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000000111?????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?00?000?11???????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111110001010?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110100?0?11???????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010000?0?11???????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111111010010?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?00111101000010?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110100001010????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111?0??11??1111?????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111100100111?????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111110110111?????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010010111?????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111?1011011?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011111001?011?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001111010?1011?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?0011110101?011?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    26'b0?001110000??011?1????????  :  v_ldst_dest_incr[7] = 1'b1;
	    default : v_ldst_dest_incr[7] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b0?00111000001010?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111000110?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111110000111?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111001111?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111010001?0001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111101000001?0001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111000111?0001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100010?0?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?1000000?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100?1010?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?1010010?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110?0000?0011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?000000?0001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?001001?0001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111100?000?0001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000000?1??011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?0011??011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111101010011??001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000001???001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001100??011??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010110?0?011??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000?011??001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?????0011101000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000101010011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100001?0?0?011??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?100??011??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000110???011??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100001?00??011??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100100?1??011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b000011111?0?????0011101000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?1011011??011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110110?1??011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b00001111?10?????0011101000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010010?1??011?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000001?1??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?011011??001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001001???001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?0111??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111101101???001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110100101???001?0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?1011000??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111100011010011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001?000??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010?1000??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111000011110011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111100111110011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100011?1??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110101?00??011??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000??000??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111101000110001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000?11???11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110100000110001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111100011110001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111000000?0????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100010?010011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?100000010011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100?101010011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?101001010011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111001001?0????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110?000010011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?0?1110??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?00000010001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100??110??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?0?0101??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?101011???11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?00100110001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?100?101??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111100?00010001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111000000011??????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?101?111??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110??101??11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110100?11???11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000000?11?011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?00111?011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010100111?001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000001?1?001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111101000010?0????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001100?1011??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010110?01011??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000?0111?001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111110010011??????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100001?0?01011??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?100?1011??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111011011??????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000110??1011??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b000011111?0?111?10110?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?01?11???11??0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100001?00?1011??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100100?11?011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111101001011??????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?10110111?011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110110?11?011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010010?11?011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000001?1?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000001?11?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?0110111?001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001001?1?001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?01111?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111101101?1?001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110100101?1?001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?1011000?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?10110001?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001?000?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010?1000?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001?0001?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010?10001?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110101?000?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?10110?1?1011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100011?1?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000??000?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100011?11?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110101?00?1011??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001?0?1?1011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000??0001?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010?10?1?1011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110101?0?1?1011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?101101??1001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000?0?11?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000?11??111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000??0?1?1011?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011100000?11?1?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001?01??1001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010?101??1001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110101?01??1001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111100000010????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000??01??1001?????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?0?1110?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111100100110????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?0?11101?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100??110?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?0?0101?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?101011??111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100??1101?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?0?01011?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?101011?1?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?100?101?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?100?1011?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110??101?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000000111?????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?101?1111?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110??1011?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110100?11??111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110100?11?1?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010??111?111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110100001010????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111100100111?????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?01?11??111??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111110110111?????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111?01?11?1?11??????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010010111?????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111?1011011?1????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011111001?011?1????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001111010?1011?1????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?0011110101?011?1????????  :  v_ldst_dest_incr[6] = 1'b1;
	    26'b0?001110000??011?1????????  :  v_ldst_dest_incr[6] = 1'b1;
	    default : v_ldst_dest_incr[6] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b0?00111111010001?0001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111101000001?0001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111000001010?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111000111?0001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?000000?0001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?001001?0001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111100?000?0001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111000110?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001100??01?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110000111?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010110?0?01?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111001111?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111101010011??001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000001???001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?0?0?01?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?100??01?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000110???01?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001100??011??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010110?0?011??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?011??001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?00??01?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?????0011101000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?0?0?011??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000001?1??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?100??011??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000110???011??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?00??011??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b000011111?0?????0011101000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?0111??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b00001111?10?????0011101000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100?1010?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110?0000?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000001?1??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?011011??001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001001???001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?0111??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111101101???001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?1011000??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100101???001?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100010?0?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?000??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?1000000?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?1000??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?1010010?001??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?1011000??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100011?1??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?00??01?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??000??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000000?1??01??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?000??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?1000??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?0011??01??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100011?1??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?00??011??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?11???1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??000??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111101000110001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?11???11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100000110001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000010101001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111100011110001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?1110??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111000000?0????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100100?1??01??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?1011011??01??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110110?1??01??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100??110??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010010?1??01??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?0101??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101011???1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111001001?0????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?1110??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?100?101??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?00000010001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101?111??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110??101??1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100??110??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?0101??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100?11???1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101011???11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?00100110001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?100?101??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111100?00010001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111000000011??????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101?111??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110??101??11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100?11???11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110001101001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001100?101?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100001111001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010110?0101?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110011111001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010100111?001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000001?1?001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?0?0101?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111101000010?0????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?100?101?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000110??101?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001100?1011??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?01?11???1?1?0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010110?01011??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?0111?001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?00?101?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000001?1?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110001001?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110010011??????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?0?01011??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000001?11?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110001001?10?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?100?1011??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111011011??????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000110??1011??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b000011111?0?111?10110?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?01?11???11??0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111010001?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100001?00?1011??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111101001011??????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?01111?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111010001?10?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111101000001?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000001?1?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111101000001?10?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100?10101001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110?00001001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000001?11?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0110111?001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001001?1?001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?01111?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111101101?1?001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?10110001?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100101?1?001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100010?01001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?0001?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?10000001001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?10001?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?1011000?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?10100101001??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?10110001?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??000?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100011?11?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?00?101?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?000?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??0001?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000000?11?01??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?1000?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?0001?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?10001?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?000?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?00111?01??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?0?11?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100011?1?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?11??11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??000?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100011?11?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?00?1011??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?11?1?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??0001?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111000110?1?1??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101101??1001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000?0?11?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?11??111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110000111?11???????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011100000?11?1?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?01??1001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110000111?1?1??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?101??1001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111001111?1?1??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?01??1001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?01?000?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111000110?11???????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?11101?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111100000010????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??01??1001?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100100?11?01??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?10110111?01??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110110?11?01??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?0101?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101011??11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100??1101?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010010?11?01??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?01011?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111001111?11???????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?1110?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010??000?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?00?101?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101011?1?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?100?101?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111100100110????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?11101?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?100?1011?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101?111?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110??101?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100??110?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?0101?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100010?0?11???????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101?1111?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110??1011?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100?11??11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101011??111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100??1101?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0?01011?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100010?0?1?1??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100?11?1?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101011?1?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?100?101?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?100?1011?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110??101?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110100?0?1?1??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000000111?????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?101?1111?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110??1011?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010000?0?1?1??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100?11??111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100?11?1?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010??111?111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?10110?1?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111110001010?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110100?0?11???????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010000?0?11???????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111111010010?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?0?1?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?0??110?11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?10?1?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?00111101000010?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?0?1?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110100001010????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?01?11?1?1?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??0?1?101??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100??11??11?1?????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111100100111?????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?01?11??111??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111110110111?????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111?01?11?1?11??????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010010111?????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111?1011011?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011111001?011?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001111010?1011?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?0011110101?011?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    26'b0?001110000??011?1????????  :  v_ldst_dest_incr[5] = 1'b1;
	    default : v_ldst_dest_incr[5] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b010011111?0?111?00100?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111010001?0001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111101000001?0001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111000001010?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111000111?0001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?000000?0001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?001001?0001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111100?000?0001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111000110?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111110000111?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111001111?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111101010011??001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100000001???001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100000?011??001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?????0011101000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b000011111?0?????0011101000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b00001111?10?????0011101000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100?1010?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110?0000?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?011011??001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001001???001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111101101???001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110100101???001?0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100010?0?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?1000000?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?1010010?001??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000000?1??01??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?0011??01??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111101000110001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110100000110001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000010101001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111100011110001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111000000?0????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100100?1??01??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001100??01???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010110?0?01???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?1011011??01??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110110?1??01??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010010?1??01??0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111001001?0????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100001?0?0?01???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?100??01???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000110???01???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100001?00??01???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?00000010001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000001?1??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?00100110001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111100?00010001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?0111??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111000000011??????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110001101001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100001111001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110011111001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?1011000??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010100111?001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100000001?1?001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001?000??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111101000010?0????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010?1000??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100000?0111?001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100011?1??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110101?00??01???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000??000??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111110010011??????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111011011??????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b000011111?0?111?10110?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111101001011??????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100000?11???1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100?10101001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110?00001001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?0110111?001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001001?1?001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111101101?1?001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110100101?1?001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100010?01001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?10000001001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?0?1110??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?10100101001??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100??110??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?0?0101??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000000?11?01??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?101011???1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?00111?01??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?100?101??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?101?111??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110??101??1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110100?11???1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?101101??1001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001?01??1001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010?101??1001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110101?01??1001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111100000010????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000??01??1001?????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100100?11?01??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001100?101???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010110?0101???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?10110111?01??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110110?11?01??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010010?11?01??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111100100110????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100001?0?0101???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?100?101???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000110??101???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?01?11???1???0000  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100001?00?101???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000001?1?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000001?11?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?01111?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000000111?????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?10110?1?101??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?1011000?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?10110001?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001?0?1?101??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010?10?1?101??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001?000?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010?1000?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110101?0?1?101??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001?0001?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110100001010????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010?10001?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110101?000?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100011?1?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000??0?1?101??????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000??000?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100011?11?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110101?00?101???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000??0001?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100100111?????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110110111?????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000?0?11?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010010111?????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100000?11??11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011100000?11?1?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?0?1110?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?0?11101?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100??110?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?0?0101?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?101011??11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111100??1101?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?1011011?1????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?0?01011?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?101011?1?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?100?101?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?100?1011?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111001?011?1????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110??101?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010?1011?1????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111?101?1111?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111110??1011?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110100?11??11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110101?011?1????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011110100?11?1?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001111010??111?11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?001110000??011?1????????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?01?11??11???????  :  v_ldst_dest_incr[4] = 1'b1;
	    26'b0?0011111?01?11?1?1???????  :  v_ldst_dest_incr[4] = 1'b1;
	    default : v_ldst_dest_incr[4] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b010011111?0?111?00100?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111000001010?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111000110?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111110000111?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111001111?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?????00?1101000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111000000??1??011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110?0000?00?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?0?11??011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010000?0?00?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?000111?00?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b000011111?0?????00?1101000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100011??00?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b00001111?10?????00?1101000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100?1010?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110?0000?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100?111?00?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000000?1??0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?0011??0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100010?0?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?1000000?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101?00???011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?1010010?001??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00?000?00?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000000?1??01??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?0011??01??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000??1???011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100100?1??0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110110?1??0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111000111?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101001???0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010010?1??0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000010101001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?1011??0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000?01???0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100100?1??01??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001100??01???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111010001?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010110?0?01???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?1011011??01??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110110?1??01??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0??11???011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010010?1??01??0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?000000?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100001?0?0?01???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?100??01???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?0101???11?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?0????011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000110???01???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111101000001?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?10????011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100001?00??01???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00?101???11?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?100?101???11?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100?000?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101?111???11?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??0????011?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110??101???11?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?011????11?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?01101???0?1?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000001?1??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100?11????11?0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?0111??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110001101001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111101010011??????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000001???????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100001111001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110011111001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?1011000??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?001001?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000?011??????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?000??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111101000010?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?1000??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111000000??1?1011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100011?1??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101?00??01???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111000000??11?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110?0000100?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??000??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?0?111?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010000?0100?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b000011111?0?111?10110?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?000111100?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100011?100?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000?11???1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?011011??????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100?10101001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111101101???????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110?00001001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100?111100?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000000?11?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?00111?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100010?01001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10000001001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?1110??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101?00?1?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001001???????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10100101001??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100011??1??1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00?000100?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100??110??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100101???????0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?0101??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000000?11?01??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101011???1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?000111?1??1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?00111?01??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000??1?1?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?100?101??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100?111?1??1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101?111??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110??101??1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?0?11?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100?11???1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100100?11?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111000110?1?1??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110110?11?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100011110????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111110000111?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101001?1?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010010?11?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111110000111?1?1??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111001111?1?1??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?10111?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111000110?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000?01?1?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100100?11?01??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001100?101???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111101000110????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010110?0101???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10110111?01??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110110?11?01??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00100??1??1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0??11?1?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110100?0?1??1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010010?11?01??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111001111?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00000010????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?01?1?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111010001?1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010000?0?1??1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100001?0?0101???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?100?101???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?01011??11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?0??1?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000110??101???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00?1?1?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100000110????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111101000001?1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?10??1?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?01?11???1???0000  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?100?1?1?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111000111?1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100001?00?101???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00?1011??11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100010?0?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?100?1011??11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100?00010????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??0???1011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110??1?1?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10?011??1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000??1??1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100010?0?1?1??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000001?1?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10110?1?10?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101?1111??11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??0??1?011?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110??1011??11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?011?1??11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?01101?1?0?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?100?11??1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111110001001?1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000001?11?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100?11?1??11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110100?0?1?1??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10??111?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?0?1?10?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?01111?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?10?1?10?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010000?0?1?1??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101?0?1?10?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??0?1?10?1?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10110?1?101??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010100111?????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111110001010?1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000001?1?????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110100?0?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?1011000?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?10110001?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010000?0?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111111010010?1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?0?1?101??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?00100110????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111000000??1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?10?1?101??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?000?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000?0111?????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111100100??1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?00111101000010?1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?1000?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101?0?1?101??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?0001?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?01?0?0?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100001010????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?10001?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101?000?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100011?1?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??0?1?101??????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??000?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100011?11?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101?00?101???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??0001?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010??0?0?1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000?0?11?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000?11??11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011100000?11?1?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0110111?????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111101101?1?????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?1110?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?11101?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001001?1?????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100??110?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?0101?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101011??11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111100??1101?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100101?1?????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0?01011?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101011?1?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?100?101?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?0??11??1?11?????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?100?1011?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110??101?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101?1111?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111110??1011?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100?11??11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110100?11?1?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010??111?11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111?101101??1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111001?01??1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001111010?101??1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011110101?01??1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?01?11??11???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?0011111?01?11?1?1???????  :  v_ldst_dest_incr[3] = 1'b1;
	    26'b0?001110000??01??1????????  :  v_ldst_dest_incr[3] = 1'b1;
	    default : v_ldst_dest_incr[3] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b010011111?0?111?00100?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?????00?1101000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110?0000?00?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010000?0?00?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?000111?00?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b000011111?0?????00?1101000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111100011??00?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b00001111?10?????00?1101000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111100?111?00?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000000?1??0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?0011??0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100010?0?001??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?1000000?001??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?1010010?001??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?00?000?00?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111000000??1??01??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?0?11??01??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100100?1??0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110110?1??0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111111000111?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101001???0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010010?1??0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?1011??0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000?01???0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001100??01???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111111010001?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010110?0?01???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?000000?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100001?0?0?01???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?100??01???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101?00??001??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000110???01???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111101000001?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100001?00??01???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111100?000?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?01101???0?1?0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000001?1??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000??1???01??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?0111??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111101010011??????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000001???????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?1011000??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?001001?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000?011??????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?000??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111101000010?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?1000??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100011?1??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101?00??01???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0??11??001??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110?0000100?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??000??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010000?0100?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?0101???1??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?0????01??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b000011111?0?111?10110?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?000111100?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?10????01??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?00?101???1??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111100011?100?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?100?101???1??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000?11???1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?011011??????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111101101???????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101?111???1??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??0????01??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110??101???1??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?011????1??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111100?111100?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100?11????1??0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000000?11?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?00111?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100010?01001??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?10000001001??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?1110??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001001???????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?10100101001??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?00?000100?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100??110??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100101???????0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?0101??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101011???1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?100?101??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111000000??1?101??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101?111??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110??101??1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?00111000000??11?01??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100?11???1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?0?111?01??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100100?11?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110110?11?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111100011110????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101001?1?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010010?11?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?10111?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000?01?1?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001100?101???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111101000110????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010110?0101???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?00000010????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100001?0?0101???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?100?101???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101?00?1001??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?1001110?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000110??101???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100000110????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?01?11???1???0000  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100001?00?101???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111100?00010????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000001?1?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?10110?1?10?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?01101?1?0?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000001?11?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000??1?1?01??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?0?1?10?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?01111?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?10?1?10?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?0?11?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101?0?1?10?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??0?1?10?1?????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010100111?????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000001?1?????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?1011000?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?10110001?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?00100110????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?000?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000?0111?????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?1000?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?0001?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100001010????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?10001?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101?000?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100011?1?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?10110???101??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??000?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100011?11?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101?00?101???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0??11?1001??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??0001?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100??110?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?0???101??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0101?1?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100?111??1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?10???101??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?01011??1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?0??1?01??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?00?101?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000?0?11?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?10??1?01??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101?0???101??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?100?101?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000?11??11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?00?1011??1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?100?1011??1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000?11?1?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0110111?????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??0???101??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110??101?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?011??1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011100000??1??1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111101101?1?????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101?1111??1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??0??1?01??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110??1011??1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?011?1??1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100?11?1??1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010??111?1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?1110?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?11101?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001001?1?????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100??110?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?0101?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101011??11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111100??1101?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100101?1?????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?0?01011?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101011?1?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?100?101?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?100?1011?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110??101?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?01?11??1?1??????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101?1111?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111110??1011?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100?11??11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110100?11?1?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010??111?11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111?101101??1????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111001?01??1????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001111010?101??1????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011110101?01??1????????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?01?11??11???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?0011111?01?11?1?1???????  :  v_ldst_dest_incr[2] = 1'b1;
	    26'b0?001110000??01??1????????  :  v_ldst_dest_incr[2] = 1'b1;
	    default : v_ldst_dest_incr[2] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b0?001110000?????000?101000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b000011111?0?????000?101000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b00001111?10?????000?101000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?????0011101000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b000011111?0?????0011101000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b00001111?10?????0011101000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111000000??1??01??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0?11??01??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110?0000?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001100??01???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111111010001?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?000111?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010110?0?01???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111100011??0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010000?0?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100001?0?0?01???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?100??01???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?00??001??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000110???01???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111100?111?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111101000001?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111000000??1????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100001?00??01???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0?11????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000000?1??????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0011??????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000001?1??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000??1???01??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0111??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?000?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?1011000??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?001001?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?00?????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?01?1?0??1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?10?011??0??1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?000??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100100?1??????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?1000??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?101????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?11??0??1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?1?1?0??1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110110?1??????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010010?1??????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100011?1??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??1?1?0??1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110101?00??01???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0??11??001??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??000??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?1011??????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000??1?????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110101001???????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?0101???1??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?0????01??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000?01???????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?10????01??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010??111????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?101???1??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?101???1??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000?11???1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?111???1??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0????01??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??101???1??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?011????1??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100?11????1??0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?1110??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001001???????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0??11??0??1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01101???????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100??110??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100101???????0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?0101??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?0??????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101011???1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?10??????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?101??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111000000??1?101??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?111??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??101??1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0??????1?0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111000000??11?01??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100?11???1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0?111?01??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110?000010????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111111000110?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001100?101???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111101000110????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00011110????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010110?0101???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111100011?10????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010000?010????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111110000111?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111111001111?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100001?0?0101???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111000000??1?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?100?101???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?00?1001??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?1001110?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000110??101???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111100?11110????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100000110????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01?11???1???0000  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111000000??11???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100001?00?101???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0?11?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0?111???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000000?11?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000001?1?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?00111?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?00111110001001?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000001?11?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000??1?1?01??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?01111?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0?11?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100010?0?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?1011000?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?00010????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110100?0?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?10110001?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010000?0?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00100110????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0101?1?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?000?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?00?1???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?01?110??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?1000?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?10?011?10??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?101?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?0001?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100100?11?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?101?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?10001?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110101?000?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?1011???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?11?10??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?1?110??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110110?11?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100011?1?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?10110???101??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?011??1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111101?1?1?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??000?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010010?11?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100011?11?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??1?110??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110101?00?101???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000??1??1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0??11?1001??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100?11??1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0001?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?10111?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000??1?1???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100??110?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?0???101??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0101?1?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100?111??1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110101001?1?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?10???101??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010??111?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?01011??1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?0??1?01??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000?01?1?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?101?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000?0?11?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?10??1?01??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110101?0???101??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010??1111???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?101?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000?11??11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?00?1011??1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?1011??1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000?11?1?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0???101??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??101?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?011??1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011100000??1??1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?1111??1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0??1?01??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??1011??1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?011?1??1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100?11?1??1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010??111?1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01?0?0?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?1110?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0??110?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?111??1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01?001?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?11101?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001001?1?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0??11?10??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100??110?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?0101?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01101?1?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010??0?0?1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101011??11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111100??1101?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100101?1?????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?0?01011?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010??001?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?0??1???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101011?1?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?10??1???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?101?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0?1?1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?100?1011?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??101?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0???1??1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01?11??1?1??????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101?1111?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111110??1011?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??0??1???1?????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100?11??11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110100?11?1?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010??111?11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111?101101??1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111001?01??1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001111010?101??1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011110101?01??1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01?11??11???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?0011111?01?11?1?1???????  :  v_ldst_dest_incr[1] = 1'b1;
	    26'b0?001110000??01??1????????  :  v_ldst_dest_incr[1] = 1'b1;
	    default : v_ldst_dest_incr[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[5], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[1], mop[0], nf[2], nf[1], nf[0], SrcB[4], SrcB[3], SrcB[2], SrcB[1], SrcB[0]})
	    26'b0?001110000?????0000?01000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b000011111?0?????0000?01000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b00001111?10?????0000?01000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b00001111110??01100001?0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001110000?????00?1101000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b000011111?0?????00?1101000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b00001111?10?????00?1101000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010000?0?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?00111101000001?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?00111000000??1??????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?00?000?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001110000?0?11??????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?001001?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011110101001???????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?00111110001010?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?101?00??0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?0?01?1?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?10?011??0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?00111111010010?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?00?101??????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?100?11??0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?100?1?1?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?00111110000001?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111110??1?1?0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011100000??1???????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010??111??????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?01101???????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?0??11??0????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111001?0????????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010?10????????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001110000??0????????0000  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010000?010????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011110100000110????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?00111000000??1?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?00111000000??11?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001110000?0?11?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?00?00010????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001110000?0?111?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?00100110????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?0?1110?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011110101001?1?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111100??110?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?0101?1?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111000101010????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111100?111??1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?101?00?10????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?0?01?110????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?101011??1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?10?011?10????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?00?101?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?100?101?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111101001010????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?00?1011?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?100?11?10????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?100?1?110????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111000000110????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111101?1?1?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111110??1?110????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011100000??1??1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011110100?11??1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011100000??1?1?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010??111?1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010??1111?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?01101?1?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111?10110???1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111?0??11?10????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111001?0???1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010?10???1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011111001?0??1?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001111010?10??1?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?0011110101?0???1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001110000??0???1????????  :  v_ldst_dest_incr[0] = 1'b1;
	    26'b0?001110000??0??1?????????  :  v_ldst_dest_incr[0] = 1'b1;
	    default : v_ldst_dest_incr[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_ldst_index_incr (
input [6:0] Opcode,
input [2:0] funct3,
input [2:0] sew,
input [2:0] lmul,
input [1:0] mop,
input [2:0] nf,
output reg [7:0] v_ldst_index_incr
);

always_comb begin
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001110000100111  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011111?0010001  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011111000?0001  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011111000100?1  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011110101?0111  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011100000101?1  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011111001101?1  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011110101001?1  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001110000000101  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001110000000011  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111110001111  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111110110101  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111100100101  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111010010101  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_incr[7] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011111?0100011  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011110100?0011  :  v_ldst_index_incr[7] = 1'b1;
	    16'b00011110100000?1  :  v_ldst_index_incr[7] = 1'b1;
	    default : v_ldst_index_incr[7] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001110000000101  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001110000000011  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001110000000111  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110001111  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110110101  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111100100101  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111010010101  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111100010?01  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110110111  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111100100111  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111010010111  :  v_ldst_index_incr[6] = 1'b1;
	    16'b00011111?0100011  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111110100101  :  v_ldst_index_incr[6] = 1'b1;
	    16'b00011110100?0011  :  v_ldst_index_incr[6] = 1'b1;
	    16'b0001111010000101  :  v_ldst_index_incr[6] = 1'b1;
	    16'b00011110100000?1  :  v_ldst_index_incr[6] = 1'b1;
	    16'b00011111000?0011  :  v_ldst_index_incr[6] = 1'b1;
	    16'b00011111?0000001  :  v_ldst_index_incr[6] = 1'b1;
	    16'b00011111100100?1  :  v_ldst_index_incr[6] = 1'b1;
	    default : v_ldst_index_incr[6] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b00011100000101?1  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011111001101?1  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011110101001?1  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001110000000101  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001110000000011  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001110000000111  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110001111  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110110101  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111100100101  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111010010101  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111100010?01  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110110111  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111100100111  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111010010111  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011111?0100011  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111110100101  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011110100?0011  :  v_ldst_index_incr[5] = 1'b1;
	    16'b0001111010000101  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011110100000?1  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011111000?0011  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011111?0000001  :  v_ldst_index_incr[5] = 1'b1;
	    16'b00011111100100?1  :  v_ldst_index_incr[5] = 1'b1;
	    default : v_ldst_index_incr[5] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001110000000101  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001110000000011  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001110000000111  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110001111  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110110101  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111100100101  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111010010101  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111100010?01  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110110111  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111100100111  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111010010111  :  v_ldst_index_incr[4] = 1'b1;
	    16'b00011111?0100011  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111110100101  :  v_ldst_index_incr[4] = 1'b1;
	    16'b00011110100?0011  :  v_ldst_index_incr[4] = 1'b1;
	    16'b0001111010000101  :  v_ldst_index_incr[4] = 1'b1;
	    16'b00011110100000?1  :  v_ldst_index_incr[4] = 1'b1;
	    16'b00011111000?0011  :  v_ldst_index_incr[4] = 1'b1;
	    16'b00011111?0000001  :  v_ldst_index_incr[4] = 1'b1;
	    16'b00011111100100?1  :  v_ldst_index_incr[4] = 1'b1;
	    default : v_ldst_index_incr[4] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001110000100111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111100?00011  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111?10010011  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111?10000001  :  v_ldst_index_incr[3] = 1'b1;
	    16'b00011110101?0111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b00011100000101?1  :  v_ldst_index_incr[3] = 1'b1;
	    16'b00011111001101?1  :  v_ldst_index_incr[3] = 1'b1;
	    16'b00011110101001?1  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001110000000011  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001110000000111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111100010?01  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111110110111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111100100111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111010010111  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111110100101  :  v_ldst_index_incr[3] = 1'b1;
	    16'b0001111010000101  :  v_ldst_index_incr[3] = 1'b1;
	    default : v_ldst_index_incr[3] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001110000000101  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001110000000011  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001110000000111  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110001111  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110110101  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111100100101  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111010010101  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111100010?01  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110110111  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111100100111  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111010010111  :  v_ldst_index_incr[2] = 1'b1;
	    16'b00011111?0100011  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111110100101  :  v_ldst_index_incr[2] = 1'b1;
	    16'b00011110100?0011  :  v_ldst_index_incr[2] = 1'b1;
	    16'b0001111010000101  :  v_ldst_index_incr[2] = 1'b1;
	    16'b00011110100000?1  :  v_ldst_index_incr[2] = 1'b1;
	    16'b00011111000?0011  :  v_ldst_index_incr[2] = 1'b1;
	    16'b00011111?0000001  :  v_ldst_index_incr[2] = 1'b1;
	    16'b00011111100100?1  :  v_ldst_index_incr[2] = 1'b1;
	    default : v_ldst_index_incr[2] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001111100?10101  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111110100011  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111010000011  :  v_ldst_index_incr[1] = 1'b1;
	    16'b00011100000101?1  :  v_ldst_index_incr[1] = 1'b1;
	    16'b00011111001101?1  :  v_ldst_index_incr[1] = 1'b1;
	    16'b00011110101001?1  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001110000000101  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001110000000111  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111110001111  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111110110101  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111100100101  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111010010101  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111110110111  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111100100111  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111010010111  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111110100101  :  v_ldst_index_incr[1] = 1'b1;
	    16'b0001111010000101  :  v_ldst_index_incr[1] = 1'b1;
	    16'b00011111000?0011  :  v_ldst_index_incr[1] = 1'b1;
	    16'b00011111?0000001  :  v_ldst_index_incr[1] = 1'b1;
	    16'b00011111100100?1  :  v_ldst_index_incr[1] = 1'b1;
	    default : v_ldst_index_incr[1] = 1'b0;
	endcase
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001110000000101  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001110000000011  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001110000000111  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110001111  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110110101  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111100100101  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111010010101  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111100010?01  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110110111  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111100100111  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111010010111  :  v_ldst_index_incr[0] = 1'b1;
	    16'b00011111?0100011  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111110100101  :  v_ldst_index_incr[0] = 1'b1;
	    16'b00011110100?0011  :  v_ldst_index_incr[0] = 1'b1;
	    16'b0001111010000101  :  v_ldst_index_incr[0] = 1'b1;
	    16'b00011110100000?1  :  v_ldst_index_incr[0] = 1'b1;
	    16'b00011111000?0011  :  v_ldst_index_incr[0] = 1'b1;
	    16'b00011111?0000001  :  v_ldst_index_incr[0] = 1'b1;
	    16'b00011111100100?1  :  v_ldst_index_incr[0] = 1'b1;
	    default : v_ldst_index_incr[0] = 1'b0;
	endcase
end
endmodule

module autogen_v_ldst_index_reset (
input [6:0] Opcode,
input [2:0] funct3,
input [2:0] sew,
input [2:0] lmul,
input [1:0] mop,
input [2:0] nf,
output reg [7:0] v_ldst_index_reset
);

always_comb begin
	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0], nf[2], nf[1], nf[0]})
	    19'b00011100000?01?1001  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001110000000?11011  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111?10100101001  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011110100?0101001  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?0100011011  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111110?10011011  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111?10010011011  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?0001111?11  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111100?1111?11  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111100011?1?11  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?01?0101001  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?001001101?  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?00100110?1  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111110?00001?11  :  v_ldst_index_reset[7] = 1'b1;
	    19'b000111111010001101?  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111?10000001?11  :  v_ldst_index_reset[7] = 1'b1;
	    19'b000111101000001101?  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111101000110?1  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011110100000110?1  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111110001111?1?  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111110001111??1  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?00?0001?11  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001110000?00111???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111100111111??  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?00011111??  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011100000?0111???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111100011011??  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?0000001?1?  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111100?0001?1?  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?0000001??1  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111100?0001??1  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111101000011??  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011110100000011??  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111100010101???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111110100101???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111010000101???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111?10110111???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011110101?0111???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111010?10111???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111001?0111???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111100000011???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111110010011???  :  v_ldst_index_reset[7] = 1'b1;
	    19'b00011111?00?00011??  :  v_ldst_index_reset[7] = 1'b1;
	    19'b0001111110000001???  :  v_ldst_index_reset[7] = 1'b1;
	    default : v_ldst_index_reset[7] = 1'b0;
	endcase
v_ldst_index_reset[6] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_ldst_index_reset[6]

	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0], nf[2], nf[1]})
	    18'b000111000000001101  :  v_ldst_index_reset[5] = 1'b1;
	    18'b000111110010001101  :  v_ldst_index_reset[5] = 1'b1;
	    18'b000111111011001101  :  v_ldst_index_reset[5] = 1'b1;
	    18'b000111101001001101  :  v_ldst_index_reset[5] = 1'b1;
	    18'b00011111000011111?  :  v_ldst_index_reset[5] = 1'b1;
	    18'b0001111100001111?1  :  v_ldst_index_reset[5] = 1'b1;
	    18'b0001111110011111?1  :  v_ldst_index_reset[5] = 1'b1;
	    18'b0001111110001101?1  :  v_ldst_index_reset[5] = 1'b1;
	    18'b00011111000100011?  :  v_ldst_index_reset[5] = 1'b1;
	    18'b00011111100111111?  :  v_ldst_index_reset[5] = 1'b1;
	    18'b0001111100010001?1  :  v_ldst_index_reset[5] = 1'b1;
	    18'b00011111100011011?  :  v_ldst_index_reset[5] = 1'b1;
	    18'b0001111110100001?1  :  v_ldst_index_reset[5] = 1'b1;
	    18'b0001111010000001?1  :  v_ldst_index_reset[5] = 1'b1;
	    18'b00011111101000011?  :  v_ldst_index_reset[5] = 1'b1;
	    18'b00011110100000011?  :  v_ldst_index_reset[5] = 1'b1;
	    default : v_ldst_index_reset[5] = 1'b0;
	endcase
v_ldst_index_reset[4] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_ldst_index_reset[4]

	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0], nf[2], nf[1], nf[0]})
	    19'b00011100000000110?1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b000111000000001101?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b000111110010001101?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b000111111011001101?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b000111101001001101?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111000011111??  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111100001111?1?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111110011111?1?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111?01000110?1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111101?00110?1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111110001101?1?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111000100011??  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011110100?00110?1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011100000?0101???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111100111111??  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111100010001?1?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111100011011??  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111010100101???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111110100001?1?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111010000001?1?  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111?0001111??1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111100?1111??1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111100011?1??1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111010010101???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111101000011??  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111110001111???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011110100000011??  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111?0010001??1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111101000?1??1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011110100000?1??1  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111?0110101???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111100010011???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b00011111001?0101???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111110100011???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111100000001???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111010000011???  :  v_ldst_index_reset[3] = 1'b1;
	    19'b0001111110010001???  :  v_ldst_index_reset[3] = 1'b1;
	    default : v_ldst_index_reset[3] = 1'b0;
	endcase
v_ldst_index_reset[2] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_ldst_index_reset[2]

	casez({Opcode[6], Opcode[4], Opcode[3], Opcode[2], Opcode[1], Opcode[0], funct3[2], funct3[1], funct3[0], sew[2], sew[1], sew[0], lmul[2], lmul[1], lmul[0], mop[0]})
	    16'b0001110000000011  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111100001111  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111110011111  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111110001101  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111100100011  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111110110011  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111100010001  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111010010011  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111110100001  :  v_ldst_index_reset[1] = 1'b1;
	    16'b0001111010000001  :  v_ldst_index_reset[1] = 1'b1;
	    default : v_ldst_index_reset[1] = 1'b0;
	endcase
v_ldst_index_reset[0] = 1'b0; // Assigning Default value of 0
// No logic driving this. Skipping Output for v_ldst_index_reset[0]

end
endmodule

//spyglass enable_block OneModule-ML
//spyglass enable_block W398
